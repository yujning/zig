// 
// Copyright (c) 2014-2024 by SHENZHEN PANGO MICROSYSTEMS CO.,LTD
// ALL RIGHTS RESERVED.
// 
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
// 

module GTP_ADC_E2
#(
    parameter [15:0] CREG_00H = 16'h0001,
    parameter [15:0] CREG_01H = 16'hC83F,
    parameter [15:0] CREG_02H = 16'h0009,
    parameter [13:0] CREG_31H = 14'h0000,
    parameter [15:0] CREG_03H = 16'h0000,
    parameter [15:0] CREG_04H = 16'h0000,
    parameter [15:0] CREG_0AH = 16'h0000,
    parameter [15:0] CREG_05H = 16'h0000,
    parameter [15:0] CREG_06H = 16'h0000,
    parameter [15:0] CREG_0CH = 16'h0000,
    parameter [15:0] CREG_07H = 16'h0000,
    parameter [15:0] CREG_08H = 16'h0000,
    parameter [15:0] CREG_0EH = 16'h0000,
    parameter [11:0] CREG_20H = 12'h000,
    parameter [11:0] CREG_21H = 12'h000,
    parameter [11:0] CREG_22H = 12'h000,
    parameter [11:0] CREG_23H = 12'h000,
    parameter [11:0] CREG_24H = 12'h000,
    parameter [11:0] CREG_25H = 12'h000,
    parameter [11:0] CREG_26H = 12'h000,
    parameter [11:0] CREG_27H = 12'h000,
    parameter [11:0] CREG_28H = 12'h000,
    parameter [11:0] CREG_29H = 12'h000,
    parameter [11:0] CREG_2AH = 12'hCC2,
    parameter [11:0] CREG_2BH = 12'hA5B
) (
    input [1:0] VA,
    input [31:0] VAUX,
    input DCLK,
    input [7:0] DADDR,
    input DEN,
    input SECEN,
    input DWE,
    input [15:0] DI,
    output [15:0] DO,
    output DRDY,
    input CONVST,
    input RST_N,
    input LOADSC_N,
    output OVER_TEMP,
    output LOGIC_DONE_A,
    output LOGIC_DONE_B,
    output ADC_CLK_OUT,
    output DMODIFIED,
    output [4:0] ALARM
)  ;
endmodule


module GTP_APM_E2
#(
    parameter GRS_EN = "TRUE",
    parameter integer ASYNC_RST = 0,
    parameter integer X_REG = 0,
    parameter integer XB_REG = 0,
    parameter integer Y_REG = 0,
    parameter integer Z_REG = 0,
    parameter integer P_REG = 0,
    parameter integer CXO_REG = 0,
    parameter integer CPO_REG = 0,
    parameter integer MULT_REG = 0,
    parameter integer PREADD_REG = 0,
    parameter integer MODEIN_REG = 0,
    parameter integer MODEY_REG = 0,
    parameter integer MODEZ_REG = 0,
    parameter integer X_SEL = 0,
    parameter integer XB_SEL = 0,
    parameter integer CIN_SEL = 0,
    parameter integer ROUNDMODE_SEL = 0,
    parameter integer USE_SIMD = 0,
    parameter integer USE_ACCLOW = 0,
    parameter integer USE_PREADD = 0,
    parameter integer USE_POSTADD = 0,
    parameter integer USE_MULT = 1,
    parameter [47:0] P_INIT0 = 48'h000000000000,
    parameter [47:0] P_INIT1 = 48'h000000000000
) (
    output COUT,
    output [47:0] CPO,
    output [29:0] CXO,
    output [24:0] CXBO,
    output [47:0] P,
    input CIN,
    input [47:0] CPI,
    input [29:0] CXI,
    input [24:0] CXBI,
    input [29:0] X,
    input [24:0] XB,
    input [17:0] Y,
    input [47:0] Z,
    input [4:0] MODEIN,
    input [2:0] MODEY,
    input [3:0] MODEZ,
    input CLK,
    input CEX1,
    input CEX2,
    input CEX3,
    input CEXB,
    input CEY1,
    input CEY2,
    input CEZ,
    input CEM,
    input CEP,
    input CEPRE,
    input CEMODEIN,
    input CEMODEY,
    input CEMODEZ,
    input RSTX,
    input RSTXB,
    input RSTY,
    input RSTZ,
    input RSTM,
    input RSTP,
    input RSTPRE,
    input RSTMODEIN,
    input RSTMODEY,
    input RSTMODEZ
)  ;
endmodule


module GTP_BUF
(
    output Z,
    input I
)  ;
endmodule


module GTP_CFGCLK
(
    input CLKIN,
    input CE_N
)  ;
endmodule


module GTP_CLKBUFCE
(
    output CLKOUT,
    input CE,
    input CLKIN
)  ;
endmodule


module GTP_CLKBUFG
(
    output CLKOUT,
    input CLKIN
)  ;
endmodule


module GTP_CLKBUFGCE
#(
    parameter DEFAULT_VALUE = 1'b0,
    parameter SIM_DEVICE = "TITAN"
) (
    output CLKOUT,
    input CLKIN,
    input CE
)  ;
endmodule


module GTP_CLKBUFGMUX
#(
    parameter TRIGGER_MODE = "NORMAL",
    parameter SIM_DEVICE = "TITAN"
) (
    output CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input SEL
)  ;
endmodule


module GTP_CLKBUFGMUX_E1
#(
    parameter TRIGGER_MODE = "NEGEDGE",
    parameter INIT_SEL = "CLK0"
) (
    output CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input SEL,
    input EN
)  ;
endmodule


module GTP_CLKBUFGMUX_E2
#(
    parameter TRIGGER_MODE = "NEGEDGE",
    parameter INIT_SEL = "CLK0"
) (
    output CLKOUT,
    input CLKIN0,
    input CLKIN1,
    input DETECT_CLK0,
    input DETECT_CLK1,
    input SEL
)  ;
endmodule


module GTP_CLKBUFM
(
    output CLKOUT,
    input CLKIN
)  ;
endmodule


module GTP_CLKBUFMCE
#(
    parameter CE_TYPE = "SYNC",
    parameter CE_INV = "FALSE",
    parameter TRIGGER_MODE = "POSEDGE"
) (
    output CLKOUT,
    input CLKIN,
    input CE
)  ;
endmodule


module GTP_CLKBUFR
(
    output CLKOUT,
    input CLKIN
)  ;
endmodule


module GTP_CLKBUFX
(
    output CLKOUT,
    input CLKIN
)  ;
endmodule


module GTP_CLKBUFXCE
#(
    parameter CE_TYPE = "SYNC",
    parameter CE_INV = "FALSE",
    parameter TRIGGER_MODE = "POSEDGE"
) (
    output CLKOUT,
    input CLKIN,
    input CE
)  ;
endmodule


module GTP_CLKPD
#(
    parameter CPD_EDGE = "POSEDGE",
    parameter HPIO = "FALSE"
) (
    output FLAG_PD,
    output LOCK,
    input RST,
    input CLK_SAMPLE,
    input CLK_CTRL,
    input CLK_PHY,
    input DONE
)  ;
endmodule


module GTP_DDC_E2
#(
    parameter GRS_EN = "TRUE",
    parameter CLKA_GATE_EN = "FALSE",
    parameter WCLK_DELAY_SEL = "FALSE",
    parameter DDC_MODE = "QUAD_RATE",
    parameter R_EXTEND = "FALSE",
    parameter DELAY_SEL = 1'b0,
    parameter IFIFO_GENERIC = "FALSE",
    parameter [2:0] RADDR_INIT = 3'b000,
    parameter [1:0] DATA_RATE = 2'b00
) (
    output WCLK,
    output WCLK_DELAY,
    output DQSI_DELAY,
    output DQSIB_DELAY,
    output DGTS,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    output READ_VALID,
    output [1:0] DQS_DRIFT,
    output DRIFT_DETECT_ERR,
    output DQS_DRIFT_STATUS,
    output DQS_SAMPLE,
    input RST,
    input RST_TRAINING_N,
    input CLKA,
    input CLKB,
    input DQSI,
    input DQSIB,
    input [7:0] DELAY_STEP0,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP2,
    input [7:0] DELAY_STEP3,
    input [7:0] DELAY_STEP4,
    input [3:0] DQS_GATE_CTRL,
    input GATE_SEL,
    input [1:0] CLK_GATE_CTRL,
    input CLKA_GATE
)  ;
endmodule


module GTP_DDC_E2_DFT
#(
    parameter GRS_EN = "TRUE",
    parameter DDC_MODE = "QUAD_RATE",
    parameter GATE_MODE = "DEFAULT",
    parameter CLKA_GATE_EN = "FALSE",
    parameter WCLK_DELAY_SEL = "FALSE",
    parameter R_EXTEND = "FALSE",
    parameter DELAY_SEL = 1'b0,
    parameter IFIFO_GENERIC = "FALSE",
    parameter [2:0] RADDR_INIT = 3'b000,
    parameter [1:0] DATA_RATE = 2'b00
) (
    output WCLK,
    output WCLK_DELAY,
    output DQSI_DELAY,
    output DQSIB_DELAY,
    output DGTS,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    output READ_VALID,
    output [1:0] DQS_DRIFT,
    output DRIFT_DETECT_ERR,
    output DQS_DRIFT_STATUS,
    output DQS_SAMPLE,
    output GATE_HIGHB,
    output GATE_HIGH_LATCHB,
    input RST,
    input RST_TRAINING_N,
    input CLKA,
    input CLKB,
    input DQSI,
    input DQSIB,
    input [7:0] DELAY_STEP0,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP2,
    input [7:0] DELAY_STEP3,
    input [7:0] DELAY_STEP4,
    input [3:0] DQS_GATE_CTRL,
    input GATE_SEL,
    input [1:0] CLK_GATE_CTRL,
    input CLKA_GATE
)  ;
endmodule


module GTP_DDC_E3
#(
    parameter GRS_EN = "TRUE",
    parameter DDC_MODE = "QUAD_RATE",
    parameter GATE_MODE = "DEFAULT",
    parameter CLKA_GATE_EN = "FALSE",
    parameter WCLK_DELAY_SEL = "FALSE",
    parameter R_EXTEND = "FALSE",
    parameter DELAY_SEL = 1'b0,
    parameter IFIFO_GENERIC = "FALSE",
    parameter [2:0] RADDR_INIT = 3'b000,
    parameter [1:0] DATA_RATE = 2'b00
) (
    output WCLK,
    output WCLK_DELAY,
    output DQSI_DELAY,
    output DQSIB_DELAY,
    output DGTS,
    output [2:0] IFIFO_WADDR,
    output [2:0] IFIFO_RADDR,
    output READ_VALID,
    output [1:0] DQS_DRIFT,
    output DRIFT_DETECT_ERR,
    output DQS_DRIFT_STATUS,
    output DQS_SAMPLE,
    input RST,
    input RST_TRAINING_N,
    input CLKA,
    input CLKB,
    input DQSI,
    input DQSIB,
    input [7:0] DELAY_STEP0,
    input [7:0] DELAY_STEP1,
    input [7:0] DELAY_STEP2,
    input [7:0] DELAY_STEP3,
    input [7:0] DELAY_STEP4,
    input [3:0] DQS_GATE_CTRL,
    input GATE_SEL,
    input [1:0] CLK_GATE_CTRL,
    input CLKA_GATE
)  ;
endmodule


module GTP_DFF
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK
)  ;
endmodule


module GTP_DFF_C
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK,
    input C
)  ;
endmodule


module GTP_DFF_CE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK,
    input C,
    input CE
)  ;
endmodule


module GTP_DFF_E
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK,
    input CE
)  ;
endmodule


module GTP_DFF_P
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input CLK,
    input P
)  ;
endmodule


module GTP_DFF_PE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input CLK,
    input P,
    input CE
)  ;
endmodule


module GTP_DFF_R
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK,
    input R
)  ;
endmodule


module GTP_DFF_RE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input CLK,
    input R,
    input CE
)  ;
endmodule


module GTP_DFF_S
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input CLK,
    input S
)  ;
endmodule


module GTP_DFF_SE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input CLK,
    input S,
    input CE
)  ;
endmodule


module GTP_DLATCH
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input G
)  ;
endmodule


module GTP_DLATCH_C
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input G,
    input C
)  ;
endmodule


module GTP_DLATCH_CE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input G,
    input C,
    input GE
)  ;
endmodule


module GTP_DLATCH_E
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b0
) (
    output Q,
    input D,
    input G,
    input GE
)  ;
endmodule


module GTP_DLATCH_P
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input G,
    input P
)  ;
endmodule


module GTP_DLATCH_PE
#(
    parameter GRS_EN = "TRUE",
    parameter INIT = 1'b1
) (
    output Q,
    input D,
    input G,
    input P,
    input GE
)  ;
endmodule


module GTP_DLL_E2
#(
    parameter GRS_EN = "TRUE",
    parameter [7:0] CAL_INIT = 8'b00011111,
    parameter integer DELAY_STEP_OFFSET = 0,
    parameter DELAY_SEL = 1'b0,
    parameter FAST_LOCK = "FALSE",
    parameter [1:0] FDIV = 2'b10,
    parameter INT_CLK = 1'b0,
    parameter [1:0] UPD_DLY = 2'b01,
    parameter HPIO = "FALSE"
) (
    output [7:0] DELAY_STEP,
    output [7:0] DELAY_STEP1,
    output LOCK,
    input CLKIN,
    input SYS_CLK,
    input PWD,
    input RST,
    input UPDATE_N
)  ;
endmodule


module GTP_DRM18K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter [17:0] RSTA_VAL = 18'h00000,
    parameter [17:0] RSTB_VAL = 18'h00000,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 9,
    parameter integer RAM_ADDR_WIDTH = 11,
    parameter INIT_FORMAT = "BIN"
) (
    output [17:0] DOA,
    output [17:0] DOB,
    input [17:0] DIA,
    input [17:0] DIB,
    input [13:0] ADDRA,
    input ADDRA_HOLD,
    input [13:0] ADDRB,
    input ADDRB_HOLD,
    input [3:0] BWEA,
    input [1:0] BWEB,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB
)  ;
endmodule


module GTP_DRM36K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter [2:0] CSA_MASK = 3'b000,
    parameter [2:0] CSB_MASK = 3'b000,
    parameter integer DATA_WIDTH_A = 18,
    parameter integer DATA_WIDTH_B = 18,
    parameter WRITE_MODE_A = "NORMAL_WRITE",
    parameter WRITE_MODE_B = "NORMAL_WRITE",
    parameter integer DOA_REG = 0,
    parameter integer DOB_REG = 0,
    parameter integer DOA_REG_CLKINV = 0,
    parameter integer DOB_REG_CLKINV = 0,
    parameter [35:0] RSTA_VAL = 36'h000000000,
    parameter [35:0] RSTB_VAL = 36'h000000000,
    parameter RST_TYPE = "SYNC",
    parameter RAM_MODE = "TRUE_DUAL_PORT",
    parameter RAM_CASCADE = "NONE",
    parameter ECC_READ_EN = "FALSE",
    parameter ECC_WRITE_EN = "FALSE",
    parameter [287:0] INIT_00 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_01 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_02 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_03 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_04 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_05 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_06 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_07 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_08 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_09 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_0F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_10 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_11 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_12 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_13 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_14 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_15 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_16 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_17 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_18 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_19 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_1F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_20 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_21 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_22 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_23 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_24 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_25 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_26 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_27 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_28 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_29 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_2F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_30 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_31 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_32 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_33 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_34 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_35 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_36 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_37 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_38 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_39 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_3F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_40 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_41 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_42 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_43 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_44 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_45 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_46 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_47 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_48 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_49 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_4F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_50 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_51 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_52 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_53 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_54 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_55 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_56 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_57 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_58 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_59 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_5F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_60 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_61 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_62 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_63 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_64 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_65 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_66 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_67 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_68 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_69 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_6F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_70 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_71 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_72 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_73 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_74 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_75 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_76 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_77 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_78 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_79 = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7A = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7B = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7C = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7D = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7E = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter [287:0] INIT_7F = 288'h000000000000000000000000000000000000000000000000000000000000000000000000,
    parameter INIT_FILE = "NONE",
    parameter integer BLOCK_X = 0,
    parameter integer BLOCK_Y = 0,
    parameter integer RAM_DATA_WIDTH = 18,
    parameter integer RAM_ADDR_WIDTH = 11,
    parameter INIT_FORMAT = "BIN"
) (
    output COUTA,
    output COUTB,
    output [35:0] DOA,
    output [35:0] DOB,
    output ECC_SBITERR,
    output ECC_DBITERR,
    output [8:0] ECC_RDADDR,
    output [7:0] ECC_PARITY,
    input CINA,
    input CINB,
    input [35:0] DIA,
    input [35:0] DIB,
    input [15:0] ADDRA,
    input ADDRA_HOLD,
    input [15:0] ADDRB,
    input ADDRB_HOLD,
    input [2:0] CSA,
    input [2:0] CSB,
    input [7:0] BWEA,
    input [3:0] BWEB,
    input CLKA,
    input CLKB,
    input CEA,
    input CEB,
    input WEA,
    input WEB,
    input ORCEA,
    input ORCEB,
    input RSTA,
    input RSTB,
    input INJECT_SBITERR,
    input INJECT_DBITERR
)  ;
endmodule


module GTP_EFUSECODE
#(
    parameter [31:0] SIM_EFUSE_VALUE = 32'h12345678
) (
    output [31:0] EFUSE_CODE
)  ;
endmodule


module GTP_FIFO18K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 18,
    parameter integer DO_REG = 0,
    parameter [13:0] ALMOST_FULL_OFFSET = 14'h0080,
    parameter [13:0] ALMOST_EMPTY_OFFSET = 14'h0080,
    parameter [35:0] RST_VAL = 36'h000000000,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter SYNC_FIFO = "FALSE"
) (
    output ALMOST_EMPTY,
    output ALMOST_FULL,
    output EMPTY,
    output FULL,
    output [35:0] DO,
    input [35:0] DI,
    input WCLK,
    input RCLK,
    input WCE,
    input RCE,
    input ORCE,
    input RST
)  ;
endmodule


module GTP_FIFO36K_E1
#(
    parameter GRS_EN = "TRUE",
    parameter integer DATA_WIDTH = 18,
    parameter integer DO_REG = 0,
    parameter ECC_READ_EN = "FALSE",
    parameter ECC_WRITE_EN = "FALSE",
    parameter [14:0] ALMOST_FULL_OFFSET = 15'h0080,
    parameter [14:0] ALMOST_EMPTY_OFFSET = 15'h0080,
    parameter [71:0] RST_VAL = 72'h000000000000000000,
    parameter integer USE_EMPTY = 0,
    parameter integer USE_FULL = 0,
    parameter SYNC_FIFO = "FALSE"
) (
    output ALMOST_EMPTY,
    output ALMOST_FULL,
    output EMPTY,
    output FULL,
    output [71:0] DO,
    output ECC_SBITERR,
    output ECC_DBITERR,
    input [71:0] DI,
    input WCLK,
    input RCLK,
    input WCE,
    input RCE,
    input ORCE,
    input RST,
    input INJECT_SBITERR,
    input INJECT_DBITERR
)  ;
endmodule


module GTP_GPLL
#(
    parameter real CLKIN_FREQ = 50.0,
    parameter LOCK_MODE = 1'b0,
    parameter integer STATIC_RATIOI = 1,
    parameter integer STATIC_RATIOM = 1,
    parameter real STATIC_RATIO0 = 1.0,
    parameter integer STATIC_RATIO1 = 1,
    parameter integer STATIC_RATIO2 = 1,
    parameter integer STATIC_RATIO3 = 1,
    parameter integer STATIC_RATIO4 = 1,
    parameter integer STATIC_RATIO5 = 1,
    parameter integer STATIC_RATIO6 = 1,
    parameter real STATIC_RATIOF = 1.0,
    parameter integer STATIC_DUTY0 = 2,
    parameter integer STATIC_DUTY1 = 2,
    parameter integer STATIC_DUTY2 = 2,
    parameter integer STATIC_DUTY3 = 2,
    parameter integer STATIC_DUTY4 = 2,
    parameter integer STATIC_DUTY5 = 2,
    parameter integer STATIC_DUTY6 = 2,
    parameter integer STATIC_DUTYF = 2,
    parameter integer STATIC_PHASE = 0,
    parameter integer STATIC_PHASE0 = 0,
    parameter integer STATIC_PHASE1 = 0,
    parameter integer STATIC_PHASE2 = 0,
    parameter integer STATIC_PHASE3 = 0,
    parameter integer STATIC_PHASE4 = 0,
    parameter integer STATIC_PHASE5 = 0,
    parameter integer STATIC_PHASE6 = 0,
    parameter integer STATIC_PHASEF = 0,
    parameter integer STATIC_CPHASE0 = 0,
    parameter integer STATIC_CPHASE1 = 0,
    parameter integer STATIC_CPHASE2 = 0,
    parameter integer STATIC_CPHASE3 = 0,
    parameter integer STATIC_CPHASE4 = 0,
    parameter integer STATIC_CPHASE5 = 0,
    parameter integer STATIC_CPHASE6 = 0,
    parameter integer STATIC_CPHASEF = 0,
    parameter CLK_DPS0_EN = "FALSE",
    parameter CLK_DPS1_EN = "FALSE",
    parameter CLK_DPS2_EN = "FALSE",
    parameter CLK_DPS3_EN = "FALSE",
    parameter CLK_DPS4_EN = "FALSE",
    parameter CLK_DPS5_EN = "FALSE",
    parameter CLK_DPS6_EN = "FALSE",
    parameter CLK_DPSF_EN = "FALSE",
    parameter CLK_CAS5_EN = "FALSE",
    parameter CLKOUT0_SYN_EN = "FALSE",
    parameter CLKOUT1_SYN_EN = "FALSE",
    parameter CLKOUT2_SYN_EN = "FALSE",
    parameter CLKOUT3_SYN_EN = "FALSE",
    parameter CLKOUT4_SYN_EN = "FALSE",
    parameter CLKOUT5_SYN_EN = "FALSE",
    parameter CLKOUT6_SYN_EN = "FALSE",
    parameter CLKOUTF_SYN_EN = "FALSE",
    parameter SSC_MODE = "DISABLE",
    parameter real SSC_FREQ = 50.0,
    parameter INTERNAL_FB = "CLKOUTF",
    parameter EXTERNAL_FB = "DISABLE",
    parameter BANDWIDTH = "OPTIMIZED"
) (
    output CLKOUT0,
    output CLKOUT0N,
    output CLKOUT1,
    output CLKOUT1N,
    output CLKOUT2,
    output CLKOUT2N,
    output CLKOUT3,
    output CLKOUT3N,
    output CLKOUT4,
    output CLKOUT5,
    output CLKOUT6,
    output CLKOUTF,
    output CLKOUTFN,
    output LOCK,
    output DPS_DONE,
    output [15:0] APB_RDATA,
    output APB_READY,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input DPS_CLK,
    input DPS_EN,
    input DPS_DIR,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUT5_SYN,
    input CLKOUT6_SYN,
    input CLKOUTF_SYN,
    input PLL_PWD,
    input RST,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [15:0] APB_WDATA
)  ;
endmodule


module GTP_GRS
(
    input GRS_N
)  ;
endmodule


module GTP_HPIO_VREF
#(
    parameter BANK_LOC = "BANKR5"
) (
    input [7:0] CODE_VREF0,
    input [7:0] CODE_VREF1,
    input [7:0] CODE_VREF2,
    input [7:0] CODE_VREF3
)  ;
endmodule


module GTP_HSSTHP_BUFDS
#(
    parameter PMA_CFG_COMMPOWERUP = "ON",
    parameter PMA_REG_COM_PD = "FALSE",
    parameter PMA_REG_COM_PD_OW = "FALSE",
    parameter PMA_REG_HPLL_REFCLK_PD = "ON",
    parameter PMA_REG_REFCLK_FAB = "REFCLK"
) (
    input COM_POWERDOWN,
    input PAD_REFCLKP,
    input PAD_REFCLKN,
    output REFCLK_OUTP,
    output PMA_REFCLK_TO_FABRIC
)  ;
endmodule


module GTP_HSSTHP_HPLL
#(
    parameter PMA_REG_REFCLK0_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_REFCLK1_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_PLL_JTAG0_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG0_LPF_RSEL = "20K",
    parameter PMA_REG_PLL_JTAG1_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG1_LPF_RSEL = "20K",
    parameter integer PMA_REG_IBIAS_STATIC_SEL_7_0 = 255,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_15_8 = 247,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_18_16 = 7,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_21_19 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_29_22 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_37_30 = 1,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_4_0 = 31,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_8_5 = 15,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_12_9 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_17_13 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0,
    parameter PMA_REG_CALIB_CLKDIV_RATION = "DIV1",
    parameter PMA_REG_TX_RATE_CHANGE_SEL0 = "CLK_FROM_HPLL",
    parameter PMA_REG_TX_RATE_CHANGE_SEL1 = "SEL_SYNC_RATE_CHANGE",
    parameter PMA_REG_TLING_IMPEDANCE_CTRL = "125OHM",
    parameter integer PMA_ANA_COM_REG_143 = 0,
    parameter integer PMA_ANA_COM_REG_149 = 0,
    parameter integer PMA_ANA_COM_REG_155 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_3_0 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_11_4 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_15_12 = 0,
    parameter PMA_REG_HPLL_VCOLDO_EN = "TRUE",
    parameter PMA_REG_HPLL_LDO_VOL_RANGE_O = "1000MV",
    parameter PMA_REG_HPLL_LDO_VOL_RANGE_I = "640MV",
    parameter integer PMA_REG_HPLL_REFCLK_DIV = 1,
    parameter PMA_REG_HPLL_CHARGE_PUMP_PD = "WORK",
    parameter integer PMA_REG_HPLL_CHARGE_PUMP_CTRL = 10,
    parameter PMA_REG_HPLL_VCTRL_SEL_L = "0.4V",
    parameter PMA_REG_HPLL_VCTRL_SEL_H = "0.5V",
    parameter PMA_REG_HPLL_LPF_RES_SEL = "5K",
    parameter PMA_REG_HPLL_PCURRENT_SEL = "16*IO",
    parameter integer PMA_REG_HPLL_VCO_EN = 1,
    parameter PMA_REG_HPLL_PCURRENT_SEL0 = "10*IO",
    parameter integer PMA_REG_HPLL_PCURRENT_SEL1 = 0,
    parameter integer PMA_REG_REFCLK_RST_SEL = 0,
    parameter integer PMA_REG_NFC_STIC_DIS_N = 0,
    parameter integer PMA_REG_HPLL_FBDIV0 = 20,
    parameter integer PMA_REG_HPLL_FBDIV1 = 20,
    parameter PMA_REG_HPLL_PHASE_SEL = "DIV2",
    parameter integer PMA_REG_HPLL_CFG_7_0 = 7,
    parameter integer PMA_REG_HPLL_CFG_15_8 = 132,
    parameter PMA_REG_PLL_LOCKDET_RESET_N = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_RESET_N_OW = "FALSE",
    parameter PMA_REG_READY_OR_LOCK = "FALSE",
    parameter PMA_REG_HPLL_READY = "FALSE",
    parameter PMA_REG_HPLL_READY_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_REFCT_0 = "TRUE",
    parameter integer PMA_REG_PLL_LOCKDET_REFCT_2_1 = 1,
    parameter integer PMA_REG_PLL_LOCKDET_FBCT = 3,
    parameter integer PMA_REG_PLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_REG_PLL_LOCKDET_ITER = 0,
    parameter integer PMA_REG_PLL_UNLOCKDET_ITER = 2,
    parameter PMA_REG_PLL_LOCKDET_EN_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_EN = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_MODE = "FALSE",
    parameter PMA_REG_PLL_LOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKED = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED = "FALSE",
    parameter PMA_REG_PLL_LOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_LOCKDET_REPEAT = "FALSE",
    parameter PMA_REG_NOFBCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_NOREFCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_RESCAL_EN = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_OW = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_1_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_5_2 = 0,
    parameter PMA_REG_RESCAL_I_CODE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_ITER_VALID_SEL = 0,
    parameter PMA_REG_RESCAL_WAIT_SEL = "FALSE",
    parameter integer PMA_REG_I_CTRL_MAX = 45,
    parameter integer PMA_REG_I_CTRL_MIN_1_0 = 3,
    parameter integer PMA_REG_I_CTRL_MIN_5_2 = 4,
    parameter integer PMA_REG_RESCAL_I_CODE_3_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_5_4 = 2,
    parameter PMA_REG_RESCAL_INT_R_SMALL_VAL = "FALSE",
    parameter PMA_REG_RESCAL_INT_R_SMALL_OW = "FALSE",
    parameter PMA_REG_RESCAL_I_CODE_PMA = "FALSE",
    parameter PMA_REG_REFCLK0_JTAG_OE = "FALSE",
    parameter PMA_REG_REFCLK1_JTAG_OE = "FALSE",
    parameter PMA_REG_RES_CAL_EN = "FALSE",
    parameter PMA_REG_HPLL_RSTN = "FALSE",
    parameter PMA_REG_HPLL_RSTN_OW = "FALSE",
    parameter PMA_REG_HPLL_PD = "FALSE",
    parameter PMA_REG_HPLL_PD_OW = "FALSE",
    parameter PMA_REG_LC_VCO_CAL_EN = "FALSE",
    parameter PMA_REG_DIV_CALI_BYPASS = "TRUE",
    parameter integer PMA_REG_CALIB_WAIT = 3,
    parameter integer PMA_REG_CALIB_TIMER = 0,
    parameter integer PMA_REG_BAND_LB = 0,
    parameter PMA_REG_BAND_HB_0 = "TRUE",
    parameter integer PMA_REG_BAND_HB_4_1 = 15,
    parameter PMA_CFG_HSST_RSTN = "TRUE",
    parameter PMA_CFG_PLLPOWERUP = "ON",
    parameter PMA_PLL_RSTN = "TRUE",
    parameter PMA_REG_LANE0_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE1_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE2_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE3_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_HPLL_REFCLK_SEL = "DISABLE",
    parameter integer PMA_REG_HSST_LAST_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_LAST_REFCLK1_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK1_SEL = 0,
    parameter integer PMA_ANA_COM_REG_142 = 0,
    parameter integer PMA_ANA_COM_REG_145_144 = 1,
    parameter integer PMA_ANA_COM_REG_146 = 0,
    parameter integer PMA_ANA_COM_REG_147 = 0,
    parameter integer PMA_ANA_COM_REG_148 = 0,
    parameter integer PMA_ANA_COM_REG_151_150 = 1,
    parameter integer PMA_ANA_COM_REG_152 = 0,
    parameter integer PMA_ANA_COM_REG_153 = 0,
    parameter integer PMA_ANA_COM_REG_154 = 0,
    parameter integer PMA_ANA_COM_REG_157_156 = 1,
    parameter integer PMA_ANA_COM_REG_158 = 0,
    parameter integer PMA_ANA_COM_REG_159 = 0
) (
    input P_CFG_RST_HPLL,
    input P_CFG_CLK_HPLL,
    input P_CFG_PSEL_HPLL,
    input P_CFG_ENABLE_HPLL,
    input P_CFG_WRITE_HPLL,
    input [11:0] P_CFG_ADDR_HPLL,
    input [7:0] P_CFG_WDATA_HPLL,
    output P_CFG_READY_HPLL,
    output [7:0] P_CFG_RDATA_HPLL,
    output P_CFG_INT_HPLL,
    input P_HPLL_POWERDOWN,
    input P_HPLL_RST,
    input P_HPLL_LOCKDET_RST,
    input P_RES_CAL_RST,
    input P_TX_SYNC,
    input P_HPLL_DIV_SYNC,
    input P_REFCLK_DIV_SYNC,
    input P_HPLL_VCO_CALIB_EN,
    input [5:0] P_RESCAL_I_CODE_I,
    output [5:0] P_RES_CAL_CODE_FABRIC,
    output P_HPLL_READY,
    input P_HPLL_DIV_CHANGE,
    output PMA_HPLL_READY_O,
    output PMA_HPLL_REFCLK_O,
    output PMA_TX_SYNC_HPLL_O,
    output PMA_HPLL_CK0,
    output PMA_HPLL_CK90,
    output PMA_HPLL_CK180,
    output PMA_HPLL_CK270,
    output TX_SYNC_REFSYNC_O,
    output REFCLK_SYNC_REFSYNC_O,
    output DIV_SYNC_REFSYNC_O,
    input P_HPLL_REFCLK_I,
    input REFCLK_TO_TX_SYNC_I,
    input REFCLK_TO_REFCLK_SYNC_I,
    input REFCLK_TO_DIV_SYNC_I,
    input ANA_TX_SYNC_I,
    input ANA_HPLL_REFCLK_SYNC_I,
    input ANA_HPLL_DIV_SYNC_I,
    input P_PLL_REFCLK6_I,
    input REFCLK0,
    input REFCLK1,
    input REFCLK0_FROM_UPPER_HSST,
    input REFCLK1_FROM_UPPER_HSST,
    input REFCLK0_FROM_LOWER_HSST,
    input REFCLK1_FROM_LOWER_HSST,
    input REFCLK_FROM_FABRIC,
    output LPLL_REFCKOUT_CH0,
    output LPLL_REFCKOUT_CH1,
    output LPLL_REFCKOUT_CH2,
    output LPLL_REFCKOUT_CH3,
    output REFCLK0_FOR_UPPER_HSST,
    output REFCLK1_FOR_UPPER_HSST,
    output REFCLK0_FOR_LOWER_HSST,
    output REFCLK1_FOR_LOWER_HSST,
    input TX_SYNC_FROM_UPPER_HSST,
    input TX_SYNC_FROM_LOWER_HSST,
    output TX_SYNC_FOR_UPPER_HSST,
    output TX_SYNC_FOR_LOWER_HSST,
    output ANA_TX_SYNC_O,
    input REFCLK_SYNC_FROM_UPPER_HSST,
    input REFCLK_SYNC_FROM_LOWER_HSST,
    output REFCLK_SYNC_FOR_UPPER_HSST,
    output REFCLK_SYNC_FOR_LOWER_HSST,
    input DIV_SYNC_FROM_UPPER_HSST,
    input DIV_SYNC_FROM_LOWER_HSST,
    output DIV_SYNC_FOR_UPPER_HSST,
    output DIV_SYNC_FOR_LOWER_HSST
)  ;
endmodule


module GTP_HSSTHP_HPLL_DFT
#(
    parameter PMA_REG_REFCLK0_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_REFCLK1_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_PLL_JTAG0_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG0_LPF_RSEL = "20K",
    parameter PMA_REG_PLL_JTAG1_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG1_LPF_RSEL = "20K",
    parameter integer PMA_REG_IBIAS_STATIC_SEL_7_0 = 255,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_15_8 = 247,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_18_16 = 7,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_21_19 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_29_22 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_37_30 = 1,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_4_0 = 31,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_8_5 = 15,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_12_9 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_17_13 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0,
    parameter PMA_REG_CALIB_CLKDIV_RATION = "DIV1",
    parameter PMA_REG_TX_RATE_CHANGE_SEL0 = "CLK_FROM_HPLL",
    parameter PMA_REG_TX_RATE_CHANGE_SEL1 = "SEL_SYNC_RATE_CHANGE",
    parameter PMA_REG_TLING_IMPEDANCE_CTRL = "125OHM",
    parameter integer PMA_ANA_COM_REG_143 = 0,
    parameter integer PMA_ANA_COM_REG_149 = 0,
    parameter integer PMA_ANA_COM_REG_155 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_3_0 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_11_4 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_15_12 = 0,
    parameter PMA_REG_HPLL_VCOLDO_EN = "TRUE",
    parameter PMA_REG_HPLL_LDO_VOL_RANGE_O = "1000MV",
    parameter PMA_REG_HPLL_LDO_VOL_RANGE_I = "640MV",
    parameter integer PMA_REG_HPLL_REFCLK_DIV = 1,
    parameter PMA_REG_HPLL_CHARGE_PUMP_PD = "WORK",
    parameter integer PMA_REG_HPLL_CHARGE_PUMP_CTRL = 10,
    parameter PMA_REG_HPLL_VCTRL_SEL_L = "0.4V",
    parameter PMA_REG_HPLL_VCTRL_SEL_H = "0.5V",
    parameter PMA_REG_HPLL_LPF_RES_SEL = "5K",
    parameter PMA_REG_HPLL_PCURRENT_SEL = "16*IO",
    parameter integer PMA_REG_HPLL_VCO_EN = 1,
    parameter PMA_REG_HPLL_PCURRENT_SEL0 = "10*IO",
    parameter integer PMA_REG_HPLL_PCURRENT_SEL1 = 0,
    parameter integer PMA_REG_REFCLK_RST_SEL = 0,
    parameter integer PMA_REG_NFC_STIC_DIS_N = 0,
    parameter integer PMA_REG_HPLL_FBDIV0 = 20,
    parameter integer PMA_REG_HPLL_FBDIV1 = 20,
    parameter PMA_REG_HPLL_PHASE_SEL = "DIV2",
    parameter integer PMA_REG_HPLL_CFG_7_0 = 7,
    parameter integer PMA_REG_HPLL_CFG_15_8 = 132,
    parameter PMA_REG_PLL_LOCKDET_RESET_N = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_RESET_N_OW = "FALSE",
    parameter PMA_REG_READY_OR_LOCK = "FALSE",
    parameter PMA_REG_HPLL_READY = "FALSE",
    parameter PMA_REG_HPLL_READY_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_REFCT_0 = "TRUE",
    parameter integer PMA_REG_PLL_LOCKDET_REFCT_2_1 = 1,
    parameter integer PMA_REG_PLL_LOCKDET_FBCT = 3,
    parameter integer PMA_REG_PLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_REG_PLL_LOCKDET_ITER = 0,
    parameter integer PMA_REG_PLL_UNLOCKDET_ITER = 2,
    parameter PMA_REG_PLL_LOCKDET_EN_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_EN = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_MODE = "FALSE",
    parameter PMA_REG_PLL_LOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKED = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED = "FALSE",
    parameter PMA_REG_PLL_LOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_LOCKDET_REPEAT = "FALSE",
    parameter PMA_REG_NOFBCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_NOREFCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_RESCAL_EN = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_OW = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_1_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_5_2 = 0,
    parameter PMA_REG_RESCAL_I_CODE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_ITER_VALID_SEL = 0,
    parameter PMA_REG_RESCAL_WAIT_SEL = "FALSE",
    parameter integer PMA_REG_I_CTRL_MAX = 45,
    parameter integer PMA_REG_I_CTRL_MIN_1_0 = 3,
    parameter integer PMA_REG_I_CTRL_MIN_5_2 = 4,
    parameter integer PMA_REG_RESCAL_I_CODE_3_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_5_4 = 2,
    parameter PMA_REG_RESCAL_INT_R_SMALL_VAL = "FALSE",
    parameter PMA_REG_RESCAL_INT_R_SMALL_OW = "FALSE",
    parameter PMA_REG_RESCAL_I_CODE_PMA = "FALSE",
    parameter PMA_REG_REFCLK0_JTAG_OE = "FALSE",
    parameter PMA_REG_REFCLK1_JTAG_OE = "FALSE",
    parameter PMA_REG_RES_CAL_EN = "FALSE",
    parameter PMA_REG_HPLL_RSTN = "FALSE",
    parameter PMA_REG_HPLL_RSTN_OW = "FALSE",
    parameter PMA_REG_HPLL_PD = "FALSE",
    parameter PMA_REG_HPLL_PD_OW = "FALSE",
    parameter PMA_REG_LC_VCO_CAL_EN = "FALSE",
    parameter PMA_REG_DIV_CALI_BYPASS = "TRUE",
    parameter integer PMA_REG_CALIB_WAIT = 3,
    parameter integer PMA_REG_CALIB_TIMER = 0,
    parameter integer PMA_REG_BAND_LB = 0,
    parameter PMA_REG_BAND_HB_0 = "TRUE",
    parameter integer PMA_REG_BAND_HB_4_1 = 15,
    parameter PMA_CFG_HSST_RSTN = "TRUE",
    parameter PMA_CFG_PLLPOWERUP = "ON",
    parameter PMA_PLL_RSTN = "TRUE",
    parameter PMA_REG_LANE0_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE1_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE2_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE3_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_HPLL_REFCLK_SEL = "DISABLE",
    parameter integer PMA_REG_HSST_LAST_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_LAST_REFCLK1_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK1_SEL = 0,
    parameter integer PMA_ANA_COM_REG_142 = 0,
    parameter integer PMA_ANA_COM_REG_145_144 = 1,
    parameter integer PMA_ANA_COM_REG_146 = 0,
    parameter integer PMA_ANA_COM_REG_147 = 0,
    parameter integer PMA_ANA_COM_REG_148 = 0,
    parameter integer PMA_ANA_COM_REG_151_150 = 1,
    parameter integer PMA_ANA_COM_REG_152 = 0,
    parameter integer PMA_ANA_COM_REG_153 = 0,
    parameter integer PMA_ANA_COM_REG_154 = 0,
    parameter integer PMA_ANA_COM_REG_157_156 = 1,
    parameter integer PMA_ANA_COM_REG_158 = 0,
    parameter integer PMA_ANA_COM_REG_159 = 0
) (
    input P_CFG_RST_HPLL,
    input P_CFG_CLK_HPLL,
    input P_CFG_PSEL_HPLL,
    input P_CFG_ENABLE_HPLL,
    input P_CFG_WRITE_HPLL,
    input [11:0] P_CFG_ADDR_HPLL,
    input [7:0] P_CFG_WDATA_HPLL,
    output P_CFG_READY_HPLL,
    output [7:0] P_CFG_RDATA_HPLL,
    output P_CFG_INT_HPLL,
    input P_HPLL_POWERDOWN,
    input P_HPLL_RST,
    input P_HPLL_LOCKDET_RST,
    input P_RES_CAL_RST,
    input P_TX_SYNC,
    input P_HPLL_DIV_SYNC,
    input P_REFCLK_DIV_SYNC,
    input P_HPLL_VCO_CALIB_EN,
    input [5:0] P_RESCAL_I_CODE_I,
    output [5:0] P_RES_CAL_CODE_FABRIC,
    output P_HPLL_READY,
    input P_HPLL_DIV_CHANGE,
    output PMA_HPLL_READY_O,
    output PMA_HPLL_REFCLK_O,
    output PMA_TX_SYNC_HPLL_O,
    output PMA_HPLL_CK0,
    output PMA_HPLL_CK90,
    output PMA_HPLL_CK180,
    output PMA_HPLL_CK270,
    output TX_SYNC_REFSYNC_O,
    output REFCLK_SYNC_REFSYNC_O,
    output DIV_SYNC_REFSYNC_O,
    input P_HPLL_REFCLK_I,
    input REFCLK_TO_TX_SYNC_I,
    input REFCLK_TO_REFCLK_SYNC_I,
    input REFCLK_TO_DIV_SYNC_I,
    input ANA_TX_SYNC_I,
    input ANA_HPLL_REFCLK_SYNC_I,
    input ANA_HPLL_DIV_SYNC_I,
    input P_PLL_REFCLK6_I,
    input REFCLK0,
    input REFCLK1,
    input REFCLK0_FROM_UPPER_HSST,
    input REFCLK1_FROM_UPPER_HSST,
    input REFCLK0_FROM_LOWER_HSST,
    input REFCLK1_FROM_LOWER_HSST,
    input REFCLK_FROM_FABRIC,
    output LPLL_REFCKOUT_CH0,
    output LPLL_REFCKOUT_CH1,
    output LPLL_REFCKOUT_CH2,
    output LPLL_REFCKOUT_CH3,
    output REFCLK0_FOR_UPPER_HSST,
    output REFCLK1_FOR_UPPER_HSST,
    output REFCLK0_FOR_LOWER_HSST,
    output REFCLK1_FOR_LOWER_HSST,
    input TX_SYNC_FROM_UPPER_HSST,
    input TX_SYNC_FROM_LOWER_HSST,
    output TX_SYNC_FOR_UPPER_HSST,
    output TX_SYNC_FOR_LOWER_HSST,
    output ANA_TX_SYNC_O,
    input REFCLK_SYNC_FROM_UPPER_HSST,
    input REFCLK_SYNC_FROM_LOWER_HSST,
    output REFCLK_SYNC_FOR_UPPER_HSST,
    output REFCLK_SYNC_FOR_LOWER_HSST,
    input DIV_SYNC_FROM_UPPER_HSST,
    input DIV_SYNC_FROM_LOWER_HSST,
    output DIV_SYNC_FOR_UPPER_HSST,
    output DIV_SYNC_FOR_LOWER_HSST,
    input P_TEST_SE_N,
    input P_TEST_MODE_N,
    input P_TEST_RSTN,
    input P_TEST_SI0,
    input P_TEST_SI1,
    output P_TEST_SO0,
    output P_TEST_SO1,
    input P_FOR_PMA_TEST_MODE_N,
    input P_FOR_PMA_TEST_SE_N,
    input P_FOR_PMA_TEST_CLK,
    input P_FOR_PMA_TEST_RSTN,
    input P_FOR_PMA_TEST_SI,
    output P_FOR_PMA_TEST_SO
)  ;
endmodule


module GTP_HSSTHP_HPLL_t
#(
    parameter PMA_REG_REFCLK0_FAB = "REFCLK0",
    parameter PMA_REG_REFCLK1_FAB = "REFCLK1",
    parameter integer PMA_REG_HSST_LAST_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK0_SEL = 0,
    parameter integer PMA_REG_HSST_LAST_REFCLK1_SEL = 0,
    parameter integer PMA_REG_HSST_NEXT_REFCLK1_SEL = 0,
    parameter PMA_REG_LANE0_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE1_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE2_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_LANE3_PLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_HPLL_REFCLK_SEL = "REFERENCE_CLOCK_0",
    parameter PMA_REG_REFCLK0_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_REFCLK1_IMPEDANCE_SEL = "100_OHM",
    parameter PMA_REG_PLL_JTAG0_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG0_LPF_RSEL = "20K",
    parameter PMA_REG_PLL_JTAG1_VTH_SEL = "60MV",
    parameter PMA_REG_PLL_JTAG1_LPF_RSEL = "20K",
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0,
    parameter PMA_REG_CALIB_CLKDIV_RATION = "DIV1",
    parameter PMA_REG_HPLL_REFCLK0_PD = "ON",
    parameter PMA_REG_HPLL_REFCLK1_PD = "ON",
    parameter PMA_REG_TX_RATE_CHANGE_SEL0 = "CLK_FROM_HPLL",
    parameter PMA_REG_TX_RATE_CHANGE_SEL1 = "SEL_SYNC_RATE_CHANGE",
    parameter PMA_REG_TLING_IMPEDANCE_CTRL = "125OHM",
    parameter integer PMA_ANA_COM_REG_142 = 0,
    parameter integer PMA_ANA_COM_REG_143 = 0,
    parameter integer PMA_ANA_COM_REG_145_144 = 1,
    parameter integer PMA_ANA_COM_REG_146 = 0,
    parameter integer PMA_ANA_COM_REG_147 = 0,
    parameter integer PMA_ANA_COM_REG_148 = 0,
    parameter integer PMA_ANA_COM_REG_149 = 0,
    parameter integer PMA_ANA_COM_REG_151_150 = 1,
    parameter integer PMA_ANA_COM_REG_152 = 0,
    parameter integer PMA_ANA_COM_REG_153 = 0,
    parameter integer PMA_ANA_COM_REG_154 = 0,
    parameter integer PMA_ANA_COM_REG_155 = 0,
    parameter integer PMA_ANA_COM_REG_157_156 = 1,
    parameter integer PMA_ANA_COM_REG_158 = 0,
    parameter integer PMA_ANA_COM_REG_159 = 0,
    parameter PMA_REG_COM_PD = "FALSE",
    parameter PMA_REG_COM_PD_OW = "FALSE",
    parameter integer PMA_REG_HPLL_DIV_CHANGE_3_0 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_11_4 = 0,
    parameter integer PMA_REG_HPLL_DIV_CHANGE_15_12 = 0,
    parameter PMA_REG_HPLL_VCOLDO_EN = "TRUE",
    parameter integer PMA_REG_HPLL_REFCLK_DIV = 1,
    parameter PMA_REG_HPLL_CHARGE_PUMP_PD = "WORK",
    parameter integer PMA_REG_HPLL_CHARGE_PUMP_CTRL = 10,
    parameter PMA_REG_HPLL_LPF_RES_SEL = "5K",
    parameter integer PMA_REG_HPLL_VCO_EN = 1,
    parameter integer PMA_REG_HPLL_PCURRENT_SEL1 = 0,
    parameter integer PMA_REG_REFCLK_RST_SEL = 0,
    parameter integer PMA_REG_NFC_STIC_DIS_N = 0,
    parameter integer PMA_REG_HPLL_FBDIV0 = 20,
    parameter integer PMA_REG_HPLL_FBDIV1 = 20,
    parameter PMA_REG_HPLL_PHASE_SEL = "DIV2",
    parameter integer PMA_REG_HPLL_CFG_7_0 = 7,
    parameter integer PMA_REG_HPLL_CFG_15_8 = 132,
    parameter PMA_REG_PLL_LOCKDET_RESET_N = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_RESET_N_OW = "FALSE",
    parameter PMA_REG_READY_OR_LOCK = "FALSE",
    parameter PMA_REG_HPLL_READY = "FALSE",
    parameter PMA_REG_HPLL_READY_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_REFCT_0 = "TRUE",
    parameter integer PMA_REG_PLL_LOCKDET_REFCT_2_1 = 1,
    parameter integer PMA_REG_PLL_LOCKDET_FBCT = 3,
    parameter integer PMA_REG_PLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_REG_PLL_LOCKDET_ITER = 0,
    parameter integer PMA_REG_PLL_UNLOCKDET_ITER = 2,
    parameter PMA_REG_PLL_LOCKDET_EN_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_EN = "FALSE",
    parameter PMA_REG_PLL_LOCKDET_MODE = "FALSE",
    parameter PMA_REG_PLL_LOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_LOCKED = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_OW = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED = "FALSE",
    parameter PMA_REG_PLL_LOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_PLL_UNLOCKED_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_LOCKDET_REPEAT = "FALSE",
    parameter PMA_REG_NOFBCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_NOREFCLK_STICKY_CLEAR = "FALSE",
    parameter PMA_REG_RESCAL_EN = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_OW = "FALSE",
    parameter PMA_REG_RESCAL_RST_N_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_VAL = "FALSE",
    parameter PMA_REG_RESCAL_DONE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_1_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_VAL_5_2 = 0,
    parameter PMA_REG_RESCAL_I_CODE_OW = "FALSE",
    parameter integer PMA_REG_RESCAL_ITER_VALID_SEL = 0,
    parameter PMA_REG_RESCAL_WAIT_SEL = "FALSE",
    parameter integer PMA_REG_I_CTRL_MAX = 45,
    parameter integer PMA_REG_I_CTRL_MIN_1_0 = 3,
    parameter integer PMA_REG_I_CTRL_MIN_5_2 = 4,
    parameter integer PMA_REG_RESCAL_I_CODE_3_0 = 0,
    parameter integer PMA_REG_RESCAL_I_CODE_5_4 = 2,
    parameter PMA_REG_RESCAL_INT_R_SMALL_VAL = "FALSE",
    parameter PMA_REG_RESCAL_INT_R_SMALL_OW = "FALSE",
    parameter PMA_REG_RESCAL_I_CODE_PMA = "FALSE",
    parameter PMA_REG_REFCLK0_JTAG_OE = "FALSE",
    parameter PMA_REG_REFCLK1_JTAG_OE = "FALSE",
    parameter PMA_REG_RES_CAL_EN = "FALSE",
    parameter PMA_REG_HPLL_RSTN = "FALSE",
    parameter PMA_REG_HPLL_RSTN_OW = "FALSE",
    parameter PMA_REG_HPLL_PD = "FALSE",
    parameter PMA_REG_HPLL_PD_OW = "FALSE",
    parameter PMA_REG_LC_VCO_CAL_EN = "FALSE",
    parameter PMA_REG_DIV_CALI_BYPASS = "TRUE",
    parameter integer PMA_REG_CALIB_WAIT = 3,
    parameter integer PMA_REG_CALIB_TIMER = 0,
    parameter integer PMA_REG_BAND_LB = 0,
    parameter PMA_REG_BAND_HB_0 = "TRUE",
    parameter integer PMA_REG_BAND_HB_4_1 = 15,
    parameter PMA_CFG_HSST_RSTN = "TRUE",
    parameter PMA_CFG_COMMPOWERUP = "ON",
    parameter PMA_CFG_PLLPOWERUP = "ON",
    parameter PMA_PLL_RSTN = "TRUE"
) (
    input P_CFG_RST_HPLL,
    input P_CFG_CLK_HPLL,
    input P_CFG_PSEL_HPLL,
    input P_CFG_ENABLE_HPLL,
    input P_CFG_WRITE_HPLL,
    input [11:0] P_CFG_ADDR_HPLL,
    input [7:0] P_CFG_WDATA_HPLL,
    output P_CFG_READY_HPLL,
    output [7:0] P_CFG_RDATA_HPLL,
    output P_CFG_INT_HPLL,
    input P_COM_POWERDOWN,
    input P_HPLL_POWERDOWN,
    input P_HPLL_RST,
    input P_HPLL_LOCKDET_RST,
    input P_RES_CAL_RST,
    input P_TX_SYNC,
    input P_TX_RATE_CHANGE_ON_0,
    input P_TX_RATE_CHANGE_ON_1,
    input P_HPLL_DIV_SYNC,
    input P_REFCLK_DIV_SYNC,
    input P_HPLL_VCO_CALIB_EN,
    input [5:0] P_RESCAL_I_CODE_I,
    output [5:0] P_RES_CAL_CODE_FABRIC,
    output P_REFCK2CORE_0,
    output P_REFCK2CORE_1,
    output P_HPLL_READY,
    input P_HPLL_REF_CLK,
    input P_HPLL_DIV_CHANGE,
    output PMA_HPLL_READY_LEFT,
    output PMA_HPLL_READY_RIGHT,
    output PMA_HPLL_REFCLK_LEFT,
    output PMA_HPLL_REFCLK_RIGHT,
    output PMA_LPLL_REFCKOUT_CH0,
    output PMA_LPLL_REFCKOUT_CH1,
    output PMA_LPLL_REFCKOUT_CH2,
    output PMA_LPLL_REFCKOUT_CH3,
    output [5:0] PMA_RES_CAL_LEFT,
    output [5:0] PMA_RES_CAL_RIGHT,
    output PMA_TX_RATE_CHANGE_ON0_LEFT,
    output PMA_TX_RATE_CHANGE_ON0_RIGHT,
    output PMA_TX_RATE_CHANGE_ON1_LEFT,
    output PMA_TX_RATE_CHANGE_ON1_RIGHT,
    output PMA_TX_SYNC_HPLL_LEFT,
    output PMA_TX_SYNC_HPLL_RIGHT,
    output PMA_TX_SYNC_LEFT,
    output PMA_TX_SYNC_RIGHT,
    output PMA_HPLL_CK0_CH0,
    output PMA_HPLL_CK0_CH1,
    output PMA_HPLL_CK0_CH2,
    output PMA_HPLL_CK0_CH3,
    output PMA_HPLL_CK90_CH0,
    output PMA_HPLL_CK90_CH1,
    output PMA_HPLL_CK90_CH2,
    output PMA_HPLL_CK90_CH3,
    output PMA_HPLL_CK180_CH0,
    output PMA_HPLL_CK180_CH1,
    output PMA_HPLL_CK180_CH2,
    output PMA_HPLL_CK180_CH3,
    output PMA_HPLL_CK270_CH0,
    output PMA_HPLL_CK270_CH1,
    output PMA_HPLL_CK270_CH2,
    output PMA_HPLL_CK270_CH3,
    inout [7:0] PMA_IPN50U_IN,
    input [10:0] P_FROM_LOWER_HSST_BUS,
    input [10:0] P_FROM_UPPER_HSST_BUS,
    output [10:0] P_FOR_LOWER_HSST_BUS,
    output [10:0] P_FOR_UPPER_HSST_BUS,
    input PAD_REFCLKN_0,
    input PAD_REFCLKP_0,
    input PAD_REFCLKN_1,
    input PAD_REFCLKP_1
)  ;
endmodule


module GTP_HSSTHP_LANE
#(
    parameter PCS_DYN_DLY_SEL_RX = "FALSE",
    parameter PCS_PMA_RCLK_POLINV = "PMA_RCLK",
    parameter PCS_PCS_RCLK_SEL = "RCLK",
    parameter PCS_GEAR_RCLK_SEL = "RCLK",
    parameter PCS_RCLK2FABRIC_SEL = "HARD_1",
    parameter PCS_SCAN_INTERVAL_RX = "4_CLOCKS",
    parameter PCS_BRIDGE_RCLK_SEL = "RCLK",
    parameter PCS_RCLK_POLINV = "RCLK",
    parameter PCS_TO_FABRIC_CLK_SEL = "PMA_RCLK",
    parameter PCS_CLK2ALIGNER_SEL = "TO_FABRIC_CLK",
    parameter PCS_TO_FABRIC_CLK_DIV_EN = "FALSE",
    parameter PCS_AUTO_NEAR_LOOP_EN = "FALSE",
    parameter PCS_PCS_RCLK_EN = "FALSE",
    parameter PCS_BRIDGE_PCS_RCLK_EN_SEL = "HARD_1",
    parameter PCS_BRIDGE_RCLK_EN_SEL = "HARD_0",
    parameter PCS_GEAR_RCLK_EN_SEL = "HARD_0",
    parameter PCS_NEGEDGE_EN_RX = "FALSE",
    parameter PCS_PCS_RX_RSTN = "FALSE",
    parameter PCS_BRIDGE_PCS_RSTN = "FALSE",
    parameter PCS_TO_FABRIC_RST_EN = "FALSE",
    parameter PCS_BYPASS_GEAR_RRSTN = "FALSE",
    parameter PCS_BYPASS_BRIDGE_RRSTN = "FALSE",
    parameter PCS_ALIGNER_EN_RX = "FALSE",
    parameter PCS_RX_SLAVE = "MASTER",
    parameter integer PCS_RX_CA = 0,
    parameter integer PCS_SUM_THRESHOLD_RX = 0,
    parameter integer PCS_AVG_CYCLES_RX = 0,
    parameter PCS_REG_PMA_RX2TX_PLOOP_EN = "FALSE",
    parameter PCS_REG_PMA_RX2TX_PLOOP_FIFOEN = "FALSE",
    parameter integer PCS_STEP_SIZE_RX = 0,
    parameter integer PCS_REV_CNT_LIMIT_RX = 0,
    parameter integer PCS_FILTER_CNT_SIZE_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_3_0 = 0,
    parameter integer PCS_DLY_REC_SIZE_RX = 0,
    parameter integer PCS_ALIGN_THRD_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_4 = 0,
    parameter PCS_CFG_DEC_TYPE_EN = "FALSE",
    parameter PCS_RXBRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_GE_AUTO_EN = "FALSE",
    parameter PCS_RXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_RXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_IFG_EN = "FALSE",
    parameter PCS_FLP_FULL_CHK_EN = "FALSE",
    parameter PCS_FLP_EMPTY_CHK_EN = "FALSE",
    parameter PCS_RX_POLARITY_INV = "DELAY",
    parameter PCS_FARLP_PWR_REDUCTION = "FALSE",
    parameter PCS_RXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_WDALIGN_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXDEC_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXTEST_PWR_REDUCTION = "NORMAL",
    parameter integer PCS_WA_SOS_DET_TOL = 0,
    parameter integer PCS_WA_SE_DET_TOL = 0,
    parameter PCS_RX_SAMPLE_UNION = "FALSE",
    parameter PCS_NEAR_LOOP = "FALSE",
    parameter PCS_BYPASS_WORD_ALIGN = "FALSE",
    parameter PCS_BYPASS_DENC = "FALSE",
    parameter PCS_RX_ERRCNT_CLR = "FALSE",
    parameter PCS_RX_CODE_MODE = "DUAL_8B10B",
    parameter PCS_RX_BYPASS_GEAR = "FALSE",
    parameter PCS_ERRDETECT_SILENCE = "FALSE",
    parameter PCS_RX_DATA_MODE = "8BIT",
    parameter PCS_CA_DYN_CLY_EN_RX = "FALSE",
    parameter PCS_CFG_APATTERN_STATUS_DELAY = "DELAY_ONE_CYCLE",
    parameter PCS_RX_PRBS_MODE = "DISABLE",
    parameter PCS_ALIGN_MODE = "1GB",
    parameter PCS_COMMA_DET_MODE = "PATTERN_DETECT",
    parameter integer PCS_RAPID_VMIN_1 = 0,
    parameter integer PCS_RAPID_VMIN_2 = 0,
    parameter PCS_RXBU_WIDER_EN = "40/20BIT",
    parameter integer PCS_RAPID_IMAX = 0,
    parameter PCS_RX_SPLIT = "SPLIT_22BIT_11BIT",
    parameter integer PCS_RXBRG_END_PACKET_9_8 = 0,
    parameter integer PCS_RXBRG_END_PACKET_7_0 = 0,
    parameter integer PCS_CTC_MAX_DEL = 0,
    parameter integer PCS_COMMA_REG0_9_8 = 0,
    parameter integer PCS_COMMA_REG1_9_8 = 0,
    parameter integer PCS_COMMA_MASK_9_8 = 0,
    parameter integer PCS_COMMA_REG0_7_0 = 0,
    parameter integer PCS_COMMA_REG1_7_0 = 0,
    parameter integer PCS_COMMA_MASK_7_0 = 0,
    parameter integer PCS_FLP_WRADDR_START = 0,
    parameter integer PCS_FLP_RDADDR_START = 0,
    parameter PCS_CFG_RX_BRIDGE_CLK_POLINV = "FALSE",
    parameter PCS_CTC_MODE_RD_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AFULL = 0,
    parameter PCS_FAST_LOCK_GEAR_EN = "FALSE",
    parameter PCS_CTC_MODE_WR_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AEMPTY = 0,
    parameter PCS_CTC_MODE = "ONE_BYTE",
    parameter PCS_RXBRIDGE_MODE = "BYPASS",
    parameter integer PCS_CTC_ADD_MAX = 0,
    parameter PCS_CFG_PHDET_EN_RX = "FALSE",
    parameter integer PCS_WA_SDS_DET_TOL = 0,
    parameter PCS_CEB_MODE = "10GB",
    parameter PCS_APATTERN_MODE = "ONE_BYTE",
    parameter PCS_A_REG0_8 = "FALSE",
    parameter integer PCS_RXBRG_WADDR_START = 0,
    parameter PCS_A_REG1_8 = "FALSE",
    parameter integer PCS_RXBRG_RADDR_START = 0,
    parameter integer PCS_A_REG0_7_0 = 0,
    parameter integer PCS_A_REG1_7_0 = 0,
    parameter integer PCS_CEB_RAPIDLS_MMAX = 0,
    parameter integer PCS_CEB_DETECT_TIME = 0,
    parameter integer PCS_WL_FIFO_RD = 0,
    parameter integer PCS_SKIP_REG0_9_8 = 0,
    parameter integer PCS_SKIP_REG0_7_0 = 0,
    parameter integer PCS_CFG_CONTI_SKP_SET = 0,
    parameter PCS_CFG_RX_BASE_ADV_MODE = "BASE_MODE",
    parameter integer PCS_SKIP_REG1_9_8 = 0,
    parameter integer PCS_SKIP_REG2_9_8 = 0,
    parameter integer PCS_SKIP_REG3_9_8 = 0,
    parameter integer PCS_SKIP_REG1_7_0 = 0,
    parameter integer PCS_SKIP_REG2_7_0 = 0,
    parameter integer PCS_SKIP_REG3_7_0 = 0,
    parameter integer PCS_CFG_PRBS_ERR_O_SEL = 0,
    parameter integer PCS_CFG_PD_DELAY_RX = 0,
    parameter integer PCS_WR_START_GAP = 0,
    parameter integer PCS_MIN_IFG = 0,
    parameter PCS_INT_RX_MASK_0 = "FALSE",
    parameter PCS_INT_RX_MASK_1 = "FALSE",
    parameter PCS_INT_RX_MASK_2 = "FALSE",
    parameter PCS_INT_RX_MASK_3 = "FALSE",
    parameter PCS_INT_RX_MASK_4 = "FALSE",
    parameter PCS_INT_RX_MASK_5 = "FALSE",
    parameter PCS_INT_RX_CLR_5 = "FALSE",
    parameter PCS_INT_RX_CLR_4 = "FALSE",
    parameter PCS_INT_RX_CLR_3 = "FALSE",
    parameter PCS_INT_RX_CLR_2 = "FALSE",
    parameter PCS_INT_RX_CLR_1 = "FALSE",
    parameter PCS_INT_RX_CLR_0 = "FALSE",
    parameter PCS_EM_CNT_RD_EN = "FALSE",
    parameter PCS_EM_CTRL_SEL = "SIGNAL_CTRL",
    parameter PCS_EM_MODE_CTRL = "HOLD",
    parameter PCS_EM_RD_CONDITION = "TRIGGER",
    parameter integer PCS_EM_SP_PATTERN_7_0 = 0,
    parameter integer PCS_EM_SP_PATTERN_15_8 = 0,
    parameter integer PCS_EM_SP_PATTERN_23_16 = 0,
    parameter integer PCS_EM_SP_PATTERN_31_24 = 0,
    parameter integer PCS_EM_SP_PATTERN_39_32 = 0,
    parameter integer PCS_EM_SP_PATTERN_47_40 = 0,
    parameter integer PCS_EM_SP_PATTERN_55_48 = 0,
    parameter integer PCS_EM_SP_PATTERN_63_56 = 0,
    parameter integer PCS_EM_SP_PATTERN_71_64 = 0,
    parameter integer PCS_EM_SP_PATTERN_79_72 = 0,
    parameter integer PCS_EM_PMA_MASK_7_0 = 0,
    parameter integer PCS_EM_PMA_MASK_15_8 = 0,
    parameter integer PCS_EM_PMA_MASK_23_16 = 0,
    parameter integer PCS_EM_PMA_MASK_31_24 = 0,
    parameter integer PCS_EM_PMA_MASK_39_32 = 0,
    parameter integer PCS_EM_PMA_MASK_47_40 = 0,
    parameter integer PCS_EM_PMA_MASK_55_48 = 0,
    parameter integer PCS_EM_PMA_MASK_63_56 = 0,
    parameter integer PCS_EM_PMA_MASK_71_64 = 0,
    parameter integer PCS_EM_PMA_MASK_79_72 = 0,
    parameter integer PCS_EM_EYED_MASK_7_0 = 0,
    parameter integer PCS_EM_EYED_MASK_15_8 = 0,
    parameter integer PCS_EM_EYED_MASK_23_16 = 0,
    parameter integer PCS_EM_EYED_MASK_31_24 = 0,
    parameter integer PCS_EM_EYED_MASK_39_32 = 0,
    parameter integer PCS_EM_EYED_MASK_47_40 = 0,
    parameter integer PCS_EM_EYED_MASK_55_48 = 0,
    parameter integer PCS_EM_EYED_MASK_63_56 = 0,
    parameter integer PCS_EM_EYED_MASK_71_64 = 0,
    parameter integer PCS_EM_EYED_MASK_79_72 = 0,
    parameter integer PCS_EM_PRESCALE = 0,
    parameter PCS_CFG_TEST_STATUS_SEL = "SEL_PMA_TEST_STATUS_INT",
    parameter integer PCS_CFG_DIFF_CNT_BND_RX = 0,
    parameter PCS_CFG_FLT_SEL_RX = "FALSE",
    parameter integer PCS_FILTER_BND_RX = 0,
    parameter PCS_TCLK2FABRIC_DIV_RST_M = "FALSE",
    parameter PCS_TX_PMA_TCLK_POLINV = "PMA_TCLK",
    parameter PCS_TX_TCLK_POLINV = "TCLK",
    parameter PCS_PCS_TCLK_SEL = "PMA_TCLK",
    parameter PCS_GEAR_TCLK_SEL = "PMA_TCLK",
    parameter PCS_TX_BRIDGE_TCLK_SEL = "TCLK",
    parameter PCS_TCLK2ALIGNER_SEL = "PMA_TCLK",
    parameter CA_DYN_DLY_EN_TX = "FALSE",
    parameter PCS_TX_PCS_CLK_EN_SEL = "HARDWIRED1",
    parameter PCS_TX_GEAR_CLK_EN_SEL = "HARDWIRED0",
    parameter PCS_TCLK2FABRIC_DIV_EN = "FALSE",
    parameter PCS_TCLK2FABRIC_SEL = "CLK2ALIGNER_N_DIV2",
    parameter integer DLY_ADJUST_SIZE_TX = 0,
    parameter PCS_TX_PCS_TX_RSTN = "FALSE",
    parameter PCS_TX_CA_RSTN = "FALSE",
    parameter PCS_TX_SLAVE = "MASTER",
    parameter integer PCS_TX_CA = 0,
    parameter integer PCS_CFG_PI_CLK_SEL = 0,
    parameter PCS_CFG_PI_CLK_EN_SEL = "CLK_EN_ALWAYS1",
    parameter integer PCS_CFG_PI_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_SUM_THRESHOLD_TX = 0,
    parameter integer PCS_CFG_AVG_CYCLES_TX = 0,
    parameter PCS_CFG_NEGEDGE_EN_TX = "FALSE",
    parameter integer PCS_CFG_ALIGN_THRD_TX = 0,
    parameter integer PCS_CFG_SCAN_INTERVAL_TX = 0,
    parameter integer PCS_CFG_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_REV_CNT_LIMIT_TX = 0,
    parameter integer PCS_CFG_FILTER_CNT_SIZE_TX = 0,
    parameter integer PCS_CFG_PI_DEFAULT_TX = 0,
    parameter PCS_CFG_PHDET_EN_TX = "FALSE",
    parameter PCS_PMA_TX2RX_PLOOP_EN = "FALSE",
    parameter PCS_PMA_TX2RX_SLOOP_EN = "FALSE",
    parameter PCS_CFG_DYN_DLY_SEL_TX = "FALSE",
    parameter integer PCS_CFG_DLY_REC_SIZE_TX = 0,
    parameter PCS_TX_DATA_WIDTH_MODE = "8BIT",
    parameter PCS_TX_BYPASS_BRIDGE_UINT = "FALSE",
    parameter PCS_TX_BYPASS_BRIDGE_FIFO = "FALSE",
    parameter PCS_TX_BYPASS_GEAR = "FALSE",
    parameter PCS_TX_BYPASS_ENC = "FALSE",
    parameter PCS_TX_BYPASS_BIT_SLIP = "FALSE",
    parameter PCS_TX_BRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_TXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXGEAR_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXENC_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBSLP_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_TXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_TX_ENCODER_MODE = "DUAL_8B10B",
    parameter PCS_TX_PRBS_MODE = "DISABLE",
    parameter PCS_TX_DRIVE_REG_MODE = "NO_CHANGE",
    parameter integer PCS_TX_BIT_SLIP_CYCLES = 0,
    parameter PCS_TX_BASE_ADV_MODE = "BASE",
    parameter PCS_TX_GEAR_SPLIT = "NO_SPILT",
    parameter PCS_RX_BRIDGE_CLK_POLINV = "N_CLK_INVERT",
    parameter PCS_PRBS_ERR_LPBK = "FALSE",
    parameter PCS_TX_INSERT_ER = "FALSE",
    parameter PCS_ENABLE_PRBS_GEN = "FALSE",
    parameter PCS_FAR_LOOP = "FALSE",
    parameter PCS_CFG_ENC_TYPE_EN = "FALSE",
    parameter integer PCS_TXBRG_WADDR_START = 0,
    parameter integer PCS_TXBRG_RADDR_START = 0,
    parameter PCS_CFG_TX_PIC_EN = "DISABLE",
    parameter PCS_CFG_PIC_DIRECT_INV = "FALSE",
    parameter PCS_CFG_PI_MOD_CLK_EN = "FALSE",
    parameter PCS_CFG_TX_MODULATOR_OW_EN = "FALSE",
    parameter PCS_CFG_TX_PI_SSC_MODE_EN = "FALSE",
    parameter PCS_CFG_TX_PI_OFFSET_MODE_EN = "FALSE",
    parameter integer PCS_CFG_TX_PI_SSC_MODE_SEL = 0,
    parameter PCS_CFG_TXDEEMPH_EN = "FALSE",
    parameter PCS_PI_STROBE_SEL = "FALSE",
    parameter PCS_CFG_TX_PIC_GREY_SEL = "FALSE",
    parameter PCS_CFG_PIC_RENEW_INV = "NORMAL",
    parameter integer PCS_CFG_NUM_PIC = 0,
    parameter PCS_CFG_TXPIC_OW_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_OW_VALUE_0_7 = 0,
    parameter PCS_INT_TX_MASK_0 = "FALSE",
    parameter PCS_INT_TX_MASK_1 = "FALSE",
    parameter PCS_INT_TX_MASK_2 = "FALSE",
    parameter PCS_TX_WPTR_SEL = "FALSE",
    parameter PCS_INT_TX_CLR_2 = "FALSE",
    parameter PCS_INT_TX_CLR_1 = "FALSE",
    parameter PCS_INT_TX_CLR_0 = "FALSE",
    parameter integer PCS_CFG_PD_DELAY_TX = 0,
    parameter integer PCS_CFG_DIFF_CNT_BND_TX = 0,
    parameter PCS_CFG_PD_CLK_FR_CORE_SEL = "FALSE",
    parameter PCS_CFG_FLT_SEL_TX = "FALSE",
    parameter integer PCS_FILTER_BND_TX = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_7_0 = 0,
    parameter PCS_CFG_TX_SSC_MODULATOR_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_SCALE2_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_SCALE_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_8_9 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_8 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_8_9 = 0,
    parameter PMA_REG_CHL_BIAS_POWER_SEL = "FALSE",
    parameter PMA_REG_CHL_BIAS_POWER = "FALSE",
    parameter PMA_REG_RX_BUSWIDTH = "40BIT",
    parameter PMA_REG_RX_RATE = "DIV4",
    parameter PMA_REG_RX_RATE_EN = "FALSE",
    parameter integer PMA_REG_RX_RES_TRIM = 55,
    parameter PMA_REG_RX_SIGDET_STATUS_EN = "FALSE",
    parameter integer PMA_REG_CDR_READY_THD_7_0 = 32,
    parameter integer PMA_REG_CDR_READY_THD_11_8 = 0,
    parameter PMA_REG_RX_BUSWIDTH_EN = "FALSE",
    parameter PMA_REG_RX_PCLK_EDGE_SEL = "POS_EDGE",
    parameter integer PMA_REG_RX_PIBUF_IC = 3,
    parameter integer PMA_REG_RX_DCC_IC_RX = 1,
    parameter integer PMA_REG_CDR_READY_CHECK_CTRL = 0,
    parameter PMA_REG_RX_ICTRL_TRX = "100PCT",
    parameter integer PMA_REG_PRBS_CHK_WIDTH_SEL = 1,
    parameter PMA_REG_RX_ICTRL_PIBUF = "100PCT",
    parameter PMA_REG_RX_ICTRL_PI = "100PCT",
    parameter PMA_REG_RX_ICTRL_DCC = "100PCT",
    parameter PMA_REG_TX_RATE = "DIV1",
    parameter PMA_REG_TX_RATE_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N = "TRUE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_EN = "FALSE",
    parameter PMA_REG_RX_DATA_POLARITY = "NORMAL",
    parameter PMA_REG_RX_ERR_INSERT = "FALSE",
    parameter PMA_REG_UDP_CHK_EN = "FALSE",
    parameter PMA_REG_PRBS_SEL = "PRBS7",
    parameter PMA_REG_PRBS_CHK_EN = "FALSE",
    parameter integer PMA_REG_LPLL_NFC_STIC_DIS_N = 0,
    parameter PMA_REG_BIST_CHK_PAT_SEL = "PRBS",
    parameter PMA_REG_LOAD_ERR_CNT = "FALSE",
    parameter PMA_REG_CHK_COUNTER_EN = "TRUE",
    parameter integer PMA_REG_CDR_PROP_GAN_SEL = 3,
    parameter integer PMA_REG_CDR_TUBO_PROP_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_GAIN_SEL = 2,
    parameter integer PMA_REG_CDR_TUBO_INT_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_4_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_9_5 = 28,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_2_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_9_3 = 16,
    parameter integer PMA_ANA_RX_REG_O_61_55 = 21,
    parameter integer PMA_ANA_RX_REG_O_69_62 = 0,
    parameter integer PMA_ANA_RX_REG_O_77_70 = 135,
    parameter integer PMA_ANA_RX_REG_O_85_78 = 1,
    parameter integer PMA_ANA_RX_REG_O_93_86 = 8,
    parameter integer PMA_ANA_RX_REG_O_100_94 = 64,
    parameter integer PMA_ANA_RX_REG_O_108_101 = 0,
    parameter integer PMA_ANA_RX_REG_O_111_109 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_4_0 = 3,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_5 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MAX = 11,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MIN = 15,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MAX = 35,
    parameter integer PMA_REG_COMWAKE_STATUS_CLEAR = 0,
    parameter integer PMA_REG_COMINIT_STATUS_CLEAR = 0,
    parameter PMA_REG_RX_SATA_COMINIT_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMINIT = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE = "FALSE",
    parameter PMA_REG_RX_DCC_DISABLE = "FALSE",
    parameter PMA_REG_RX_SLIP_SEL_EN = "FALSE",
    parameter integer PMA_REG_RX_SLIP_SEL_3_0 = 0,
    parameter PMA_REG_RX_SLIP_EN = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_STATUS_SEL = 5,
    parameter PMA_REG_RX_SIGDET_FSM_RST_N = "TRUE",
    parameter PMA_REG_RX_SIGDET_STATUS = "FALSE",
    parameter PMA_REG_RX_SIGDET_VTH = "36MV",
    parameter integer PMA_REG_RX_SIGDET_GRM = 0,
    parameter PMA_REG_RX_SIGDET_PULSE_EXT = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_CH2_SEL = 0,
    parameter integer PMA_REG_RX_SIGDET_CH2_CHK_WINDOW = 3,
    parameter PMA_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",
    parameter integer PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0 = 0,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3 = 0,
    parameter integer PMA_REG_RX_SIGDET_4OOB_DET_SEL = 7,
    parameter integer PMA_REG_RX_SIGDET_IC_I = 10,
    parameter integer PMA_REG_RX_EQ1_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ1_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ1_OFF = "FALSE",
    parameter integer PMA_REG_RX_EQ2_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ2_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ2_OFF = "FALSE",
    parameter integer PMA_REG_RX_ICTRL_EQ = 2,
    parameter PMA_REG_EQ_DC_CALIB_EN = "FALSE",
    parameter integer PMA_CTLE_CTRL_REG_I = 0,
    parameter PMA_CTLE_REG_FORCE_SEL_I = "FALSE",
    parameter PMA_CTLE_REG_HOLD_I = "FALSE",
    parameter integer PMA_CTLE_REG_INIT_DAC_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_INIT_DAC_I_3_2 = 0,
    parameter PMA_CTLE_REG_POLARITY_I = "FALSE",
    parameter integer PMA_CTLE_REG_SHIFTER_GAIN_I = 4,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_9_2 = 1,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_11_10 = 0,
    parameter PMA_REG_RX_RES_TRIM_EN = "FALSE",
    parameter integer PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION = 1,
    parameter integer PMA_REG_ALG_RX_TERM_VCM_SELECTION = 3,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0 = 0,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8 = 0,
    parameter PMA_REG_ALG_LOW_SPEED_MODE_ENABLE = "FALSE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER = "TRUE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION = "FALSE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_EYE_DFETAP1_PLORITY = "FALSE",
    parameter PMA_REG_CDR_SEL = "FALSE",
    parameter PMA_REG_EYE_DET_EN = "FALSE",
    parameter integer PMA_REG_PI_BIAS_CURRENT = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_6_0 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_14_7 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_21_15 = 0,
    parameter integer PMA_REG_ALG_EYE_PATH_SEL = 0,
    parameter integer PMA_REG_ALG_CTLE_TEST_SEL = 0,
    parameter PMA_REG_RX_SLIP_SEL_4 = "FALSE",
    parameter PMA_REG_ALG_RX_T1_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_CDRX_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_VP_T1_SW_PLORITY = "FALSE",
    parameter PMA_REG_ALG_RX_VP_PLORITY = "TRUE",
    parameter PMA_REG_ALG_RX_GAIN_CTRL_SUMMER = "FALSE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_T1_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_VP_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_EYE_EN = "TRUE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE = "FALSE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_REG = "FALSE",
    parameter PMA_REG_RX_PGA_OFF = "FALSE",
    parameter integer PMA_REG_ALG_CDR_XWEIGHT_I = 4,
    parameter integer PMA_REG_ALG_CDR_YWEIGHT_I = 4,
    parameter PMA_REG_ALG_CTLE_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_CTLE_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_CTLE_INITDAC_6 = 0,
    parameter PMA_REG_ALG_CTLE_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_2_0 = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_4_3 = 2,
    parameter PMA_REG_ALG_CTLEOFS_FLIPDIR_I = "TRUE",
    parameter PMA_REG_ALG_CTLEOFS_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_3_0 = 0,
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_6_4 = 4,
    parameter PMA_REG_ALG_CTLEOFS_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_SHIFT_I = 4,
    parameter PMA_REG_ALG_DFE_CTLE_PWD = "FALSE",
    parameter PMA_REG_ALG_H1_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H1_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_H1_INITDAC_6 = 0,
    parameter PMA_REG_ALG_H1_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_SHIFT_I = 4,
    parameter PMA_REG_ALG_H2_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H2_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H2_INITDAC_5_1 = 0,
    parameter PMA_REG_ALG_H2_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_SHIFT_I_1_0 = 0,
    parameter integer PMA_REG_ALG_H2_SHIFT_I_2 = 1,
    parameter PMA_REG_ALG_H3_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H3_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_INITDAC_4_0 = 0,
    parameter integer PMA_REG_ALG_H3_INITDAC_5 = 1,
    parameter PMA_REG_ALG_H3_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_SHIFT_I = 4,
    parameter PMA_REG_ALG_H4_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H4_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H4_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_H4_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_SHIFT_I = 4,
    parameter PMA_REG_ALG_H5_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H5_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_INITDAC = 16,
    parameter PMA_REG_ALG_H5_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_SHIFT_I = 4,
    parameter PMA_REG_ALG_H6_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H6_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_H6_INITDAC_4_3 = 2,
    parameter PMA_REG_ALG_H6_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_HCTLE_OFS_1_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OFS_3_2 = 2,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_6 = 1,
    parameter PMA_REG_ALG_HCTLE_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQH_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQH_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_REG_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_LEQL_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQL_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQL_REG_PRESELECT_I = 7,
    parameter integer PMA_REG_ALG_LEQL_REG_SHIFT_I = 4,
    parameter PMA_REG_ALG_NEXTBIT_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_6_0 = 127,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_14_7 = 255,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_19_15 = 31,
    parameter integer PMA_REG_ALG_SOFS_DACWIN_I = 1,
    parameter PMA_REG_ALG_SOFS_FLIP_DIR_I = "TRUE",
    parameter PMA_REG_ALG_SOFS_FORCE_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_5_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_6 = 1,
    parameter integer PMA_REG_ALG_SOFS_FORCENUM_I = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_6_3 = 8,
    parameter integer PMA_REG_ALG_SOFS_SHIFT_I = 1,
    parameter PMA_REG_ALG_SOFS_SKIP_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0 = 254,
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8 = 15,
    parameter PMA_REG_ALG_ST_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_ST_FORCEN = "FALSE",
    parameter PMA_REG_ALG_ST_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_ST_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_ST_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_ST_RECALEN = "FALSE",
    parameter integer PMA_REG_ALG_ST_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_ST_STARTCNT_7_0 = 0,
    parameter integer PMA_REG_ALG_ST_STARTCNT_15_8 = 128,
    parameter integer PMA_REG_ALG_ST_STARTCNT_19_16 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_3_0 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_11_4 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_17_12 = 2,
    parameter integer PMA_REG_ALG_ST_TOPTAP_1_0 = 3,
    parameter integer PMA_REG_ALG_ST_TOPTAP_3_2 = 3,
    parameter integer PMA_REG_ALG_SWCLK_DIV = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_3_0 = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_4 = 1,
    parameter integer PMA_REG_ALG_TAPA_NUM = 7,
    parameter integer PMA_REG_ALG_TAPB_DAC_0 = 0,
    parameter integer PMA_REG_ALG_TAPB_DAC_4_1 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_3_0 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_5_4 = 0,
    parameter integer PMA_REG_ALG_TAPC_DAC = 16,
    parameter integer PMA_REG_ALG_TAPC_NUM_0 = 1,
    parameter integer PMA_REG_ALG_TAPC_NUM_5_1 = 4,
    parameter integer PMA_REG_ALG_TAPD_DAC_2_0 = 0,
    parameter integer PMA_REG_ALG_TAPD_DAC_4_3 = 2,
    parameter integer PMA_REG_ALG_TAPD_NUM = 10,
    parameter PMA_REG_ALG_VP_FLIPDIR_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_GRN_SHIFT_I = 5,
    parameter PMA_REG_ALG_VP_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_IDEAL_2_0 = 0,
    parameter integer PMA_REG_ALG_VP_IDEAL_6_3 = 10,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_3_0 = 0,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_6_4 = 0,
    parameter PMA_REG_ALG_VP_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_VP_RED_SHIFT_I = 5,
    parameter integer PMA_REG_ALG_VPOFS_SEL_0 = 0,
    parameter integer PMA_REG_ALG_VPOFS_SEL_2_1 = 1,
    parameter integer PMA_REG_ALG_H1_UPBOUND_5_0 = 55,
    parameter integer PMA_REG_ALG_H1_UPBOUND_6 = 1,
    parameter PMA_REG_ALG_CTLEOFS_PWDN = "FALSE",
    parameter PMA_REG_ALG_LEQH_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_AGC_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_AGC_INITDAC = 10,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_1_0 = 3,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_3_2 = 0,
    parameter PMA_REG_ALG_AGC_OVERWREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_PWD = "FALSE",
    parameter integer PMA_REG_ALG_AGC_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_0 = 1,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_3_1 = 7,
    parameter integer PMA_REG_ALG_AGC_WAITSEL = 11,
    parameter PMA_REG_PI_CTRL_SEL_RX = "FALSE",
    parameter integer PMA_REG_PI_CTRL_RX_4_0 = 0,
    parameter integer PMA_REG_PI_CTRL_RX_7_5 = 0,
    parameter PMA_CFG_RX_LANE_POWERUP = "ON",
    parameter PMA_CFG_RX_PMA_RSTN = "TRUE",
    parameter PMA_INT_PMA_RX_MASK_0 = "FALSE",
    parameter PMA_INT_PMA_RX_CLR_0 = "FALSE",
    parameter PMA_CFG_CTLE_ADP_RSTN = "TRUE",
    parameter PMA_CFG_RX_CDR_RSTN = "TRUE",
    parameter PMA_CFG_RX_CLKPATH_RSTN = "TRUE",
    parameter PMA_CFG_RX_DFE_RSTN = "TRUE",
    parameter PMA_CFG_RX_LEQ_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIDING_RSTN = "TRUE",
    parameter PMA_CFG_RX_EYE_RSTN = "TRUE",
    parameter PMA_CFG_RX_CTLE_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLICER_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIP_RSTN = "TRUE",
    parameter integer PMA_REG_TX_BEACON_TIMER_SEL = 0,
    parameter PMA_REG_TX_BIT_CONV = "FALSE",
    parameter integer PMA_REG_TX_RES_CAL = 50,
    parameter integer PMA_REG_TX_UDP_DATA_20 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_26_21 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_34_27 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_39_25 = 0,
    parameter integer PMA_REG_TX_BUSWIDTH_EN = 0,
    parameter PMA_REG_TX_PD_POST = "OFF",
    parameter PMA_REG_TX_PD_POST_OW = "FALSE",
    parameter PMA_REG_TX_BUSWIDTH = "20BIT",
    parameter integer PMA_REG_EI_PCLK_DELAY_SEL = 0,
    parameter integer PMA_REG_TX_AMP_DAC0 = 25,
    parameter integer PMA_REG_TX_AMP_DAC1 = 19,
    parameter integer PMA_REG_TX_AMP_DAC2 = 14,
    parameter integer PMA_REG_TX_AMP_DAC3 = 9,
    parameter PMA_REG_TX_RXDET_THRESHOLD = "84MV",
    parameter PMA_REG_TX_BEACON_OSC_CTRL = "FALSE",
    parameter integer PMA_REG_TX_PRBS_GEN_WIDTH_SEL = 0,
    parameter PMA_REG_TX_TX2RX_SLPBACK_EN = "FALSE",
    parameter PMA_REG_TX_PCLK_EDGE_SEL = "FALSE",
    parameter PMA_REG_TX_PRBS_GEN_EN = "FALSE",
    parameter PMA_REG_TX_PRBS_SEL = "PRBS7",
    parameter integer PMA_REG_TX_UDP_DATA_7_TO_0 = 5,
    parameter integer PMA_REG_TX_UDP_DATA_15_TO_8 = 235,
    parameter integer PMA_REG_TX_UDP_DATA_19_TO_16 = 3,
    parameter integer PMA_REG_TX_FIFO_WP_CTRL = 4,
    parameter PMA_REG_TX_FIFO_EN = "FALSE",
    parameter integer PMA_REG_TX_DATA_MUX_SEL = 0,
    parameter PMA_REG_TX_ERR_INSERT = "FALSE",
    parameter PMA_REG_TX_SATA_EN = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON_OW = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON = "TRUE",
    parameter integer PMA_REG_TX_CFG_POST1 = 0,
    parameter integer PMA_REG_TX_CFG_POST2 = 0,
    parameter integer PMA_REG_TX_OOB_DELAY_SEL = 0,
    parameter PMA_REG_TX_POLARITY = "NORMAL",
    parameter PMA_REG_TX_LS_MODE_EN = "FALSE",
    parameter PMA_REG_RX_JTAG_OE = "TRUE",
    parameter integer PMA_REG_RX_ACJTAG_VHYSTSEL = 0,
    parameter PMA_REG_TX_RES_CAL_EN = "FALSE",
    parameter integer PMA_REG_RX_TERM_MODE_CTRL = 5,
    parameter PMA_REG_PLPBK_TXPCLK_EN = "FALSE",
    parameter integer PMA_REG_CLK_SEL_STROBE_TXPCLK = 2,
    parameter integer PMA_REG_TX_PH_SEL_0 = 1,
    parameter integer PMA_REG_TX_PH_SEL_6_1 = 0,
    parameter integer PMA_REG_TX_CFG_PRE = 0,
    parameter integer PMA_REG_TX_CFG_MAIN = 0,
    parameter integer PMA_REG_CFG_POST = 0,
    parameter PMA_REG_PD_MAIN = "TRUE",
    parameter PMA_REG_PD_PRE = "TRUE",
    parameter integer PMA_REG_TX_RXDET_TIMER_SEL = 87,
    parameter PMA_REG_TX_PI_CUR_BUF = "10GHz",
    parameter PMA_REG_TX_MOD_STAND_BY_EN = "FALSE",
    parameter PMA_REG_STATE_STAND_BY_SEL = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_POLAR_CTRL = "FALSE",
    parameter PMA_REG_TX_FREERUN_PD = "TRUE",
    parameter PMA_REG_TX_CHANGE_ON_SEL = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_CTRL = "FALSE",
    parameter integer PMA_REG_TX_FREERUN_RATE_0 = 0,
    parameter integer PMA_REG_TX_FREERUN_RATE_1 = 0,
    parameter PMA_REG_TX_FREERUN_RATE_OW = "FALSE",
    parameter PMA_REG_TX_RST_SYNC_CLK_SEL = "TRUE",
    parameter integer PMA_REG_TX_PI_CTRL_SEL = 0,
    parameter integer PMA_REG_TX_PI_CTRL = 0,
    parameter PMA_LANE_POWERUP = "TRUE",
    parameter PMA_POR_N = "TRUE",
    parameter PMA_TX_LANE_POWERUP = "TRUE",
    parameter PMA_TX_PMA_RSTN = "TRUE",
    parameter PMA_LPLL_POWERUP = "TRUE",
    parameter PMA_LPLL_RSTN = "TRUE",
    parameter PMA_LPLL_LOCKDET_RSTN = "TRUE",
    parameter integer PMA_REG_LPLL_PFDDELAY_SEL = 1,
    parameter PMA_REG_LPLL_PFDDELAY_EN = "TRUE",
    parameter integer PMA_REG_LPLL_VCTRL_SET = 0,
    parameter PMA_LPLL_CHARGE_PUMP_CTRL = "type",
    parameter PMA_LPLL_REFDIV = "DIV1",
    parameter integer PMA_LPLL_FBDIV = 38,
    parameter integer PMA_LPLL_LPF_RES = 1,
    parameter integer PMA_LPLL_REFLOSS_READY = 0,
    parameter integer PMA_LPLL_LOCKED_PFDDELAY = 0,
    parameter integer PMA_LPLL_MCLK_SEL = 0,
    parameter integer PMA_LPLL_TEST_SEL = 0,
    parameter PMA_LPLL_TEST_SIG_HALF_EN = "TRUE",
    parameter PMA_LPLL_TEST_V_EN = "FALSE",
    parameter PMA_LPLL_MCLK_EN = "TRUE",
    parameter integer PMA_LPLL_MCLK_DET_CTL = 16,
    parameter integer PMA_LPLL_LOCKDET_REFCT = 3,
    parameter integer PMA_LPLL_LOCKDET_FBCT = 3,
    parameter integer PMA_LPLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_LPLL_LOCKDET_ITER = 1,
    parameter integer PMA_LPLL_UNLOCKDET_ITER = 2,
    parameter integer PMA_LPLL_LOCKDET_EN_OW = 0,
    parameter integer PMA_LPLL_LOCKDET_EN = 0,
    parameter integer PMA_LPLL_LOCKDET_MODE = 0,
    parameter integer PMA_LPLL_LOCKDET_OW = 0,
    parameter integer PMA_LPLL_LOCKDETED = 0,
    parameter integer PMA_LPLL_UNLOCKDET_OW = 0,
    parameter integer PMA_LPLL_UNLOCKDETED = 0,
    parameter integer PMA_LPLL_LOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_UNLOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_LOCKDET_REPEAT = 0,
    parameter integer PMA_LPLL_NOFBCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_NOREFCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_READY_OR_LOCK = 0,
    parameter integer PMA_LPLL_READY = 0,
    parameter integer PMA_LPLL_READY_OW = 0,
    parameter PMA_REG_TXCLK_SEL = "HPLL",
    parameter PMA_REG_RXCLK_SEL = "HPLL",
    parameter integer PMA_REG_TEST_BUF = 0,
    parameter PMA_REG_RX_DEF_SEL0 = "18.75uA",
    parameter PMA_REG_RX_DEF_SEL1 = "18.75uA",
    parameter PMA_REG_TX_DIV_SEL = "25uA",
    parameter PMA_REG_LPLL_AMP_SEL = "25uA",
    parameter PMA_REG_LPLL_VCO_SEL = "25uA",
    parameter PMA_REG_LPLL_CHARGE_PUMP_SEL = "25uA",
    parameter PMA_REG_RX_EQ0_SEL = "56.25uA",
    parameter PMA_REG_RX_EQ1_SEL = "56.25uA",
    parameter PMA_REG_RX_PGA_SEL = "56.25uA",
    parameter integer PMA_REG_CHL_TEST = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_7_0 = 255,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_15_8 = 247,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_18_16 = 7,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_21_19 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_29_22 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_37_30 = 1,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_4_0 = 31,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_8_5 = 15,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_12_9 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_17_13 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0
) (
    output P_CFG_READY,
    output [7:0] P_CFG_RDATA,
    output P_CFG_INT,
    output [24:0] LANE_COUT_BUS_FORWARD,
    output [1:0] LANE_COUT_BUS_BACKWARD,
    output P_RX_PRBS_ERROR,
    output P_PCS_RX_MCB_STATUS,
    output P_PCS_LSM_SYNCED,
    output [87:0] P_RDATA,
    output P_RXDVLD,
    output P_RXDVLD_H,
    output [5:0] P_RXSTATUS,
    output [2:0] P_EM_ERROR_CNT,
    output P_LPLL_READY,
    output P_RX_SIGDET_STATUS,
    output P_RX_SATA_COMINIT,
    output P_RX_SATA_COMWAKE,
    output P_RX_LS_DATA,
    output P_RX_READY,
    output [19:0] P_TEST_STATUS,
    output P_TX_RXDET_STATUS,
    output P_RCLK2FABRIC,
    output P_TCLK2FABRIC,
    output P_CA_ALIGN_RX,
    output P_CA_ALIGN_TX,
    output P_TX_SDN,
    output P_TX_SDP,
    input P_RX_CLK_FR_CORE,
    input P_RCLK2_FR_CORE,
    input P_TX_CLK_FR_CORE,
    input P_TCLK2_FR_CORE,
    input P_PCS_RX_RST,
    input P_PCS_TX_RST,
    input P_EXT_BRIDGE_PCS_RST,
    input P_CFG_RST,
    input P_CFG_CLK,
    input P_CFG_PSEL,
    input P_CFG_ENABLE,
    input P_CFG_WRITE,
    input [11:0] P_CFG_ADDR,
    input [7:0] P_CFG_WDATA,
    input [24:0] LANE_CIN_BUS_FORWARD,
    input [1:0] LANE_CIN_BUS_BACKWARD,
    input [87:0] P_TDATA,
    input P_PCIE_EI_H,
    input P_PCIE_EI_L,
    input [15:0] P_TX_DEEMP,
    input [1:0] P_TX_DEEMP_POST_SEL,
    input P_BLK_ALIGN_CTRL,
    input P_TX_ENC_TYPE,
    input P_RX_DEC_TYPE,
    input P_PCS_BIT_SLIP,
    input P_PCS_WORD_ALIGN_EN,
    input P_RX_POLARITY_INVERT,
    input P_PCS_MCB_EXT_EN,
    input P_PCS_NEAREND_LOOP,
    input P_PCS_FAREND_LOOP,
    input P_PMA_NEAREND_PLOOP,
    input P_PMA_NEAREND_SLOOP,
    input P_PMA_FAREND_PLOOP,
    input P_PCS_PRBS_EN,
    input P_LANE_POWERDOWN,
    input P_LANE_RST,
    input P_RX_LANE_POWERDOWN,
    input P_RX_PMA_RST,
    input P_RX_CDR_RST,
    input P_RX_CLKPATH_RST,
    input P_RX_DFE_RST,
    input P_RX_LEQ_RST,
    input P_RX_SLIDING_RST,
    input P_RX_DFE_EN,
    input P_RX_T1_EN,
    input P_RX_CDRX_EN,
    input P_RX_T1_DFE_EN,
    input P_RX_T2_DFE_EN,
    input P_RX_T3_DFE_EN,
    input P_RX_T4_DFE_EN,
    input P_RX_T5_DFE_EN,
    input P_RX_T6_DFE_EN,
    input P_RX_SLIDING_EN,
    input P_RX_EYE_RST,
    input P_RX_EYE_EN,
    input [7:0] P_RX_EYE_TAP,
    input [7:0] P_RX_PIC_EYE,
    input [7:0] P_RX_PIC_FASTLOCK,
    input P_RX_PIC_FASTLOCK_STROBE,
    input P_EM_RD_TRIGGER,
    input [1:0] P_EM_MODE_CTRL,
    input P_RX_CTLE_DCCAL_RST,
    input P_RX_SLICER_DCCAL_RST,
    input P_RX_SLICER_DCCAL_EN,
    input P_RX_CTLE_DCCAL_EN,
    input P_RX_SLIP_RST,
    input P_RX_SLIP_EN,
    input P_LPLL_POWERDOWN,
    input P_LPLL_RST,
    input P_LPLL_LOCKDET_RST,
    input P_TX_LS_DATA,
    input P_TX_BEACON_EN,
    input P_TX_SWING,
    input P_TX_RXDET_REQ,
    input [1:0] P_TX_RATE,
    input [2:0] P_TX_BUSWIDTH,
    input [2:0] P_TX_FREERUN_BUSWIDTH,
    input [2:0] P_TX_MARGIN,
    input P_TX_PMA_RST,
    input P_TX_LANE_POWERDOWN,
    input P_TX_PIC_EN,
    input [1:0] P_RX_RATE,
    input [2:0] P_RX_BUSWIDTH,
    input P_RX_HIGHZ,
    input [7:0] P_CIM_CLK_ALIGNER_RX,
    input [7:0] P_CIM_CLK_ALIGNER_TX,
    input P_ALIGN_MODE_VALID_RX,
    input [1:0] P_ALIGN_MODE_RX,
    input P_ALIGN_MODE_VALID_TX,
    input [2:0] P_ALIGN_MODE_TX,
    input PMA_HPLL_CK0,
    input PMA_HPLL_CK90,
    input PMA_HPLL_CK180,
    input PMA_HPLL_CK270,
    input PMA_HPLL_READY_IN,
    input PMA_HPLL_REFCLK_IN,
    input PMA_TX_SYNC_HPLL_IN,
    input P_LPLL_REFCLK_IN,
    input P_TX_RATE_CHANGE_ON_0,
    input P_TX_RATE_CHANGE_ON_1,
    input P_TX_SYNC,
    input P_RX_SDN,
    input P_RX_SDP
)  ;
endmodule


module GTP_HSSTHP_LANE_DFT
#(
    parameter PCS_DYN_DLY_SEL_RX = "FALSE",
    parameter PCS_PMA_RCLK_POLINV = "PMA_RCLK",
    parameter PCS_PCS_RCLK_SEL = "RCLK",
    parameter PCS_GEAR_RCLK_SEL = "RCLK",
    parameter PCS_RCLK2FABRIC_SEL = "HARD_1",
    parameter PCS_SCAN_INTERVAL_RX = "4_CLOCKS",
    parameter PCS_BRIDGE_RCLK_SEL = "RCLK",
    parameter PCS_RCLK_POLINV = "RCLK",
    parameter PCS_TO_FABRIC_CLK_SEL = "PMA_RCLK",
    parameter PCS_CLK2ALIGNER_SEL = "TO_FABRIC_CLK",
    parameter PCS_TO_FABRIC_CLK_DIV_EN = "FALSE",
    parameter PCS_AUTO_NEAR_LOOP_EN = "FALSE",
    parameter PCS_PCS_RCLK_EN = "FALSE",
    parameter PCS_BRIDGE_PCS_RCLK_EN_SEL = "HARD_1",
    parameter PCS_BRIDGE_RCLK_EN_SEL = "HARD_0",
    parameter PCS_GEAR_RCLK_EN_SEL = "HARD_0",
    parameter PCS_NEGEDGE_EN_RX = "FALSE",
    parameter PCS_PCS_RX_RSTN = "FALSE",
    parameter PCS_BRIDGE_PCS_RSTN = "FALSE",
    parameter PCS_TO_FABRIC_RST_EN = "FALSE",
    parameter PCS_BYPASS_GEAR_RRSTN = "FALSE",
    parameter PCS_BYPASS_BRIDGE_RRSTN = "FALSE",
    parameter PCS_ALIGNER_EN_RX = "FALSE",
    parameter PCS_RX_SLAVE = "MASTER",
    parameter integer PCS_RX_CA = 0,
    parameter integer PCS_SUM_THRESHOLD_RX = 0,
    parameter integer PCS_AVG_CYCLES_RX = 0,
    parameter PCS_REG_PMA_RX2TX_PLOOP_EN = "FALSE",
    parameter PCS_REG_PMA_RX2TX_PLOOP_FIFOEN = "FALSE",
    parameter integer PCS_STEP_SIZE_RX = 0,
    parameter integer PCS_REV_CNT_LIMIT_RX = 0,
    parameter integer PCS_FILTER_CNT_SIZE_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_3_0 = 0,
    parameter integer PCS_DLY_REC_SIZE_RX = 0,
    parameter integer PCS_ALIGN_THRD_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_4 = 0,
    parameter PCS_CFG_DEC_TYPE_EN = "FALSE",
    parameter PCS_RXBRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_GE_AUTO_EN = "FALSE",
    parameter PCS_RXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_RXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_IFG_EN = "FALSE",
    parameter PCS_FLP_FULL_CHK_EN = "FALSE",
    parameter PCS_FLP_EMPTY_CHK_EN = "FALSE",
    parameter PCS_RX_POLARITY_INV = "DELAY",
    parameter PCS_FARLP_PWR_REDUCTION = "FALSE",
    parameter PCS_RXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_WDALIGN_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXDEC_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXTEST_PWR_REDUCTION = "NORMAL",
    parameter integer PCS_WA_SOS_DET_TOL = 0,
    parameter integer PCS_WA_SE_DET_TOL = 0,
    parameter PCS_RX_SAMPLE_UNION = "FALSE",
    parameter PCS_NEAR_LOOP = "FALSE",
    parameter PCS_BYPASS_WORD_ALIGN = "FALSE",
    parameter PCS_BYPASS_DENC = "FALSE",
    parameter PCS_RX_ERRCNT_CLR = "FALSE",
    parameter PCS_RX_CODE_MODE = "DUAL_8B10B",
    parameter PCS_RX_BYPASS_GEAR = "FALSE",
    parameter PCS_ERRDETECT_SILENCE = "FALSE",
    parameter PCS_RX_DATA_MODE = "8BIT",
    parameter PCS_CA_DYN_CLY_EN_RX = "FALSE",
    parameter PCS_CFG_APATTERN_STATUS_DELAY = "DELAY_ONE_CYCLE",
    parameter PCS_RX_PRBS_MODE = "DISABLE",
    parameter PCS_ALIGN_MODE = "1GB",
    parameter PCS_COMMA_DET_MODE = "PATTERN_DETECT",
    parameter integer PCS_RAPID_VMIN_1 = 0,
    parameter integer PCS_RAPID_VMIN_2 = 0,
    parameter PCS_RXBU_WIDER_EN = "40/20BIT",
    parameter integer PCS_RAPID_IMAX = 0,
    parameter PCS_RX_SPLIT = "SPLIT_22BIT_11BIT",
    parameter integer PCS_RXBRG_END_PACKET_9_8 = 0,
    parameter integer PCS_RXBRG_END_PACKET_7_0 = 0,
    parameter integer PCS_CTC_MAX_DEL = 0,
    parameter integer PCS_COMMA_REG0_9_8 = 0,
    parameter integer PCS_COMMA_REG1_9_8 = 0,
    parameter integer PCS_COMMA_MASK_9_8 = 0,
    parameter integer PCS_COMMA_REG0_7_0 = 0,
    parameter integer PCS_COMMA_REG1_7_0 = 0,
    parameter integer PCS_COMMA_MASK_7_0 = 0,
    parameter integer PCS_FLP_WRADDR_START = 0,
    parameter integer PCS_FLP_RDADDR_START = 0,
    parameter PCS_CFG_RX_BRIDGE_CLK_POLINV = "FALSE",
    parameter PCS_CTC_MODE_RD_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AFULL = 0,
    parameter PCS_FAST_LOCK_GEAR_EN = "FALSE",
    parameter PCS_CTC_MODE_WR_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AEMPTY = 0,
    parameter PCS_CTC_MODE = "ONE_BYTE",
    parameter PCS_RXBRIDGE_MODE = "BYPASS",
    parameter integer PCS_CTC_ADD_MAX = 0,
    parameter PCS_CFG_PHDET_EN_RX = "FALSE",
    parameter integer PCS_WA_SDS_DET_TOL = 0,
    parameter PCS_CEB_MODE = "10GB",
    parameter PCS_APATTERN_MODE = "ONE_BYTE",
    parameter PCS_A_REG0_8 = "FALSE",
    parameter integer PCS_RXBRG_WADDR_START = 0,
    parameter PCS_A_REG1_8 = "FALSE",
    parameter integer PCS_RXBRG_RADDR_START = 0,
    parameter integer PCS_A_REG0_7_0 = 0,
    parameter integer PCS_A_REG1_7_0 = 0,
    parameter integer PCS_CEB_RAPIDLS_MMAX = 0,
    parameter integer PCS_CEB_DETECT_TIME = 0,
    parameter integer PCS_WL_FIFO_RD = 0,
    parameter integer PCS_SKIP_REG0_9_8 = 0,
    parameter integer PCS_SKIP_REG0_7_0 = 0,
    parameter integer PCS_CFG_CONTI_SKP_SET = 0,
    parameter PCS_CFG_RX_BASE_ADV_MODE = "BASE_MODE",
    parameter integer PCS_SKIP_REG1_9_8 = 0,
    parameter integer PCS_SKIP_REG2_9_8 = 0,
    parameter integer PCS_SKIP_REG3_9_8 = 0,
    parameter integer PCS_SKIP_REG1_7_0 = 0,
    parameter integer PCS_SKIP_REG2_7_0 = 0,
    parameter integer PCS_SKIP_REG3_7_0 = 0,
    parameter integer PCS_CFG_PRBS_ERR_O_SEL = 0,
    parameter integer PCS_CFG_PD_DELAY_RX = 0,
    parameter integer PCS_WR_START_GAP = 0,
    parameter integer PCS_MIN_IFG = 0,
    parameter PCS_INT_RX_MASK_0 = "FALSE",
    parameter PCS_INT_RX_MASK_1 = "FALSE",
    parameter PCS_INT_RX_MASK_2 = "FALSE",
    parameter PCS_INT_RX_MASK_3 = "FALSE",
    parameter PCS_INT_RX_MASK_4 = "FALSE",
    parameter PCS_INT_RX_MASK_5 = "FALSE",
    parameter PCS_INT_RX_CLR_5 = "FALSE",
    parameter PCS_INT_RX_CLR_4 = "FALSE",
    parameter PCS_INT_RX_CLR_3 = "FALSE",
    parameter PCS_INT_RX_CLR_2 = "FALSE",
    parameter PCS_INT_RX_CLR_1 = "FALSE",
    parameter PCS_INT_RX_CLR_0 = "FALSE",
    parameter PCS_EM_CNT_RD_EN = "FALSE",
    parameter PCS_EM_CTRL_SEL = "SIGNAL_CTRL",
    parameter PCS_EM_MODE_CTRL = "HOLD",
    parameter PCS_EM_RD_CONDITION = "TRIGGER",
    parameter integer PCS_EM_SP_PATTERN_7_0 = 0,
    parameter integer PCS_EM_SP_PATTERN_15_8 = 0,
    parameter integer PCS_EM_SP_PATTERN_23_16 = 0,
    parameter integer PCS_EM_SP_PATTERN_31_24 = 0,
    parameter integer PCS_EM_SP_PATTERN_39_32 = 0,
    parameter integer PCS_EM_SP_PATTERN_47_40 = 0,
    parameter integer PCS_EM_SP_PATTERN_55_48 = 0,
    parameter integer PCS_EM_SP_PATTERN_63_56 = 0,
    parameter integer PCS_EM_SP_PATTERN_71_64 = 0,
    parameter integer PCS_EM_SP_PATTERN_79_72 = 0,
    parameter integer PCS_EM_PMA_MASK_7_0 = 0,
    parameter integer PCS_EM_PMA_MASK_15_8 = 0,
    parameter integer PCS_EM_PMA_MASK_23_16 = 0,
    parameter integer PCS_EM_PMA_MASK_31_24 = 0,
    parameter integer PCS_EM_PMA_MASK_39_32 = 0,
    parameter integer PCS_EM_PMA_MASK_47_40 = 0,
    parameter integer PCS_EM_PMA_MASK_55_48 = 0,
    parameter integer PCS_EM_PMA_MASK_63_56 = 0,
    parameter integer PCS_EM_PMA_MASK_71_64 = 0,
    parameter integer PCS_EM_PMA_MASK_79_72 = 0,
    parameter integer PCS_EM_EYED_MASK_7_0 = 0,
    parameter integer PCS_EM_EYED_MASK_15_8 = 0,
    parameter integer PCS_EM_EYED_MASK_23_16 = 0,
    parameter integer PCS_EM_EYED_MASK_31_24 = 0,
    parameter integer PCS_EM_EYED_MASK_39_32 = 0,
    parameter integer PCS_EM_EYED_MASK_47_40 = 0,
    parameter integer PCS_EM_EYED_MASK_55_48 = 0,
    parameter integer PCS_EM_EYED_MASK_63_56 = 0,
    parameter integer PCS_EM_EYED_MASK_71_64 = 0,
    parameter integer PCS_EM_EYED_MASK_79_72 = 0,
    parameter integer PCS_EM_PRESCALE = 0,
    parameter PCS_CFG_TEST_STATUS_SEL = "SEL_PMA_TEST_STATUS_INT",
    parameter integer PCS_CFG_DIFF_CNT_BND_RX = 0,
    parameter PCS_CFG_FLT_SEL_RX = "FALSE",
    parameter integer PCS_FILTER_BND_RX = 0,
    parameter PCS_TCLK2FABRIC_DIV_RST_M = "FALSE",
    parameter PCS_TX_PMA_TCLK_POLINV = "PMA_TCLK",
    parameter PCS_TX_TCLK_POLINV = "TCLK",
    parameter PCS_PCS_TCLK_SEL = "PMA_TCLK",
    parameter PCS_GEAR_TCLK_SEL = "PMA_TCLK",
    parameter PCS_TX_BRIDGE_TCLK_SEL = "TCLK",
    parameter PCS_TCLK2ALIGNER_SEL = "PMA_TCLK",
    parameter CA_DYN_DLY_EN_TX = "FALSE",
    parameter PCS_TX_PCS_CLK_EN_SEL = "HARDWIRED1",
    parameter PCS_TX_GEAR_CLK_EN_SEL = "HARDWIRED0",
    parameter PCS_TCLK2FABRIC_DIV_EN = "FALSE",
    parameter PCS_TCLK2FABRIC_SEL = "CLK2ALIGNER_N_DIV2",
    parameter integer DLY_ADJUST_SIZE_TX = 0,
    parameter PCS_TX_PCS_TX_RSTN = "FALSE",
    parameter PCS_TX_CA_RSTN = "FALSE",
    parameter PCS_TX_SLAVE = "MASTER",
    parameter integer PCS_TX_CA = 0,
    parameter integer PCS_CFG_PI_CLK_SEL = 0,
    parameter PCS_CFG_PI_CLK_EN_SEL = "CLK_EN_ALWAYS1",
    parameter integer PCS_CFG_PI_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_SUM_THRESHOLD_TX = 0,
    parameter integer PCS_CFG_AVG_CYCLES_TX = 0,
    parameter PCS_CFG_NEGEDGE_EN_TX = "FALSE",
    parameter integer PCS_CFG_ALIGN_THRD_TX = 0,
    parameter integer PCS_CFG_SCAN_INTERVAL_TX = 0,
    parameter integer PCS_CFG_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_REV_CNT_LIMIT_TX = 0,
    parameter integer PCS_CFG_FILTER_CNT_SIZE_TX = 0,
    parameter integer PCS_CFG_PI_DEFAULT_TX = 0,
    parameter PCS_CFG_PHDET_EN_TX = "FALSE",
    parameter PCS_PMA_TX2RX_PLOOP_EN = "FALSE",
    parameter PCS_PMA_TX2RX_SLOOP_EN = "FALSE",
    parameter PCS_CFG_DYN_DLY_SEL_TX = "FALSE",
    parameter integer PCS_CFG_DLY_REC_SIZE_TX = 0,
    parameter PCS_TX_DATA_WIDTH_MODE = "8BIT",
    parameter PCS_TX_BYPASS_BRIDGE_UINT = "FALSE",
    parameter PCS_TX_BYPASS_BRIDGE_FIFO = "FALSE",
    parameter PCS_TX_BYPASS_GEAR = "FALSE",
    parameter PCS_TX_BYPASS_ENC = "FALSE",
    parameter PCS_TX_BYPASS_BIT_SLIP = "FALSE",
    parameter PCS_TX_BRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_TXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXGEAR_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXENC_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBSLP_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_TXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_TX_ENCODER_MODE = "DUAL_8B10B",
    parameter PCS_TX_PRBS_MODE = "DISABLE",
    parameter PCS_TX_DRIVE_REG_MODE = "NO_CHANGE",
    parameter integer PCS_TX_BIT_SLIP_CYCLES = 0,
    parameter PCS_TX_BASE_ADV_MODE = "BASE",
    parameter PCS_TX_GEAR_SPLIT = "NO_SPILT",
    parameter PCS_RX_BRIDGE_CLK_POLINV = "N_CLK_INVERT",
    parameter PCS_PRBS_ERR_LPBK = "FALSE",
    parameter PCS_TX_INSERT_ER = "FALSE",
    parameter PCS_ENABLE_PRBS_GEN = "FALSE",
    parameter PCS_FAR_LOOP = "FALSE",
    parameter PCS_CFG_ENC_TYPE_EN = "FALSE",
    parameter integer PCS_TXBRG_WADDR_START = 0,
    parameter integer PCS_TXBRG_RADDR_START = 0,
    parameter PCS_CFG_TX_PIC_EN = "DISABLE",
    parameter PCS_CFG_PIC_DIRECT_INV = "FALSE",
    parameter PCS_CFG_PI_MOD_CLK_EN = "FALSE",
    parameter PCS_CFG_TX_MODULATOR_OW_EN = "FALSE",
    parameter PCS_CFG_TX_PI_SSC_MODE_EN = "FALSE",
    parameter PCS_CFG_TX_PI_OFFSET_MODE_EN = "FALSE",
    parameter integer PCS_CFG_TX_PI_SSC_MODE_SEL = 0,
    parameter PCS_CFG_TXDEEMPH_EN = "FALSE",
    parameter PCS_PI_STROBE_SEL = "FALSE",
    parameter PCS_CFG_TX_PIC_GREY_SEL = "FALSE",
    parameter PCS_CFG_PIC_RENEW_INV = "NORMAL",
    parameter integer PCS_CFG_NUM_PIC = 0,
    parameter PCS_CFG_TXPIC_OW_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_OW_VALUE_0_7 = 0,
    parameter PCS_INT_TX_MASK_0 = "FALSE",
    parameter PCS_INT_TX_MASK_1 = "FALSE",
    parameter PCS_INT_TX_MASK_2 = "FALSE",
    parameter PCS_TX_WPTR_SEL = "FALSE",
    parameter PCS_INT_TX_CLR_2 = "FALSE",
    parameter PCS_INT_TX_CLR_1 = "FALSE",
    parameter PCS_INT_TX_CLR_0 = "FALSE",
    parameter integer PCS_CFG_PD_DELAY_TX = 0,
    parameter integer PCS_CFG_DIFF_CNT_BND_TX = 0,
    parameter PCS_CFG_PD_CLK_FR_CORE_SEL = "FALSE",
    parameter PCS_CFG_FLT_SEL_TX = "FALSE",
    parameter integer PCS_FILTER_BND_TX = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_7_0 = 0,
    parameter PCS_CFG_TX_SSC_MODULATOR_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_SCALE2_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_SCALE_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_8_9 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_8 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_8_9 = 0,
    parameter PMA_REG_CHL_BIAS_POWER_SEL = "FALSE",
    parameter PMA_REG_CHL_BIAS_POWER = "FALSE",
    parameter PMA_REG_RX_BUSWIDTH = "40BIT",
    parameter PMA_REG_RX_RATE = "DIV4",
    parameter PMA_REG_RX_RATE_EN = "FALSE",
    parameter integer PMA_REG_RX_RES_TRIM = 55,
    parameter PMA_REG_RX_SIGDET_STATUS_EN = "FALSE",
    parameter integer PMA_REG_CDR_READY_THD_7_0 = 32,
    parameter integer PMA_REG_CDR_READY_THD_11_8 = 0,
    parameter PMA_REG_RX_BUSWIDTH_EN = "FALSE",
    parameter PMA_REG_RX_PCLK_EDGE_SEL = "POS_EDGE",
    parameter integer PMA_REG_RX_PIBUF_IC = 3,
    parameter integer PMA_REG_RX_DCC_IC_RX = 1,
    parameter integer PMA_REG_CDR_READY_CHECK_CTRL = 0,
    parameter PMA_REG_RX_ICTRL_TRX = "100PCT",
    parameter integer PMA_REG_PRBS_CHK_WIDTH_SEL = 1,
    parameter PMA_REG_RX_ICTRL_PIBUF = "100PCT",
    parameter PMA_REG_RX_ICTRL_PI = "100PCT",
    parameter PMA_REG_RX_ICTRL_DCC = "100PCT",
    parameter PMA_REG_TX_RATE = "DIV1",
    parameter PMA_REG_TX_RATE_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N = "TRUE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_EN = "FALSE",
    parameter PMA_REG_RX_DATA_POLARITY = "NORMAL",
    parameter PMA_REG_RX_ERR_INSERT = "FALSE",
    parameter PMA_REG_UDP_CHK_EN = "FALSE",
    parameter PMA_REG_PRBS_SEL = "PRBS7",
    parameter PMA_REG_PRBS_CHK_EN = "FALSE",
    parameter integer PMA_REG_LPLL_NFC_STIC_DIS_N = 0,
    parameter PMA_REG_BIST_CHK_PAT_SEL = "PRBS",
    parameter PMA_REG_LOAD_ERR_CNT = "FALSE",
    parameter PMA_REG_CHK_COUNTER_EN = "TRUE",
    parameter integer PMA_REG_CDR_PROP_GAN_SEL = 3,
    parameter integer PMA_REG_CDR_TUBO_PROP_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_GAIN_SEL = 2,
    parameter integer PMA_REG_CDR_TUBO_INT_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_4_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_9_5 = 28,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_2_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_9_3 = 16,
    parameter integer PMA_ANA_RX_REG_O_61_55 = 21,
    parameter integer PMA_ANA_RX_REG_O_69_62 = 0,
    parameter integer PMA_ANA_RX_REG_O_77_70 = 135,
    parameter integer PMA_ANA_RX_REG_O_85_78 = 1,
    parameter integer PMA_ANA_RX_REG_O_93_86 = 8,
    parameter integer PMA_ANA_RX_REG_O_100_94 = 64,
    parameter integer PMA_ANA_RX_REG_O_108_101 = 0,
    parameter integer PMA_ANA_RX_REG_O_111_109 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_4_0 = 3,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_5 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MAX = 11,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MIN = 15,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MAX = 35,
    parameter integer PMA_REG_COMWAKE_STATUS_CLEAR = 0,
    parameter integer PMA_REG_COMINIT_STATUS_CLEAR = 0,
    parameter PMA_REG_RX_SATA_COMINIT_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMINIT = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE = "FALSE",
    parameter PMA_REG_RX_DCC_DISABLE = "FALSE",
    parameter PMA_REG_RX_SLIP_SEL_EN = "FALSE",
    parameter integer PMA_REG_RX_SLIP_SEL_3_0 = 0,
    parameter PMA_REG_RX_SLIP_EN = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_STATUS_SEL = 5,
    parameter PMA_REG_RX_SIGDET_FSM_RST_N = "TRUE",
    parameter PMA_REG_RX_SIGDET_STATUS = "FALSE",
    parameter PMA_REG_RX_SIGDET_VTH = "36MV",
    parameter integer PMA_REG_RX_SIGDET_GRM = 0,
    parameter PMA_REG_RX_SIGDET_PULSE_EXT = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_CH2_SEL = 0,
    parameter integer PMA_REG_RX_SIGDET_CH2_CHK_WINDOW = 3,
    parameter PMA_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",
    parameter integer PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0 = 0,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3 = 0,
    parameter integer PMA_REG_RX_SIGDET_4OOB_DET_SEL = 7,
    parameter integer PMA_REG_RX_SIGDET_IC_I = 10,
    parameter integer PMA_REG_RX_EQ1_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ1_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ1_OFF = "FALSE",
    parameter integer PMA_REG_RX_EQ2_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ2_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ2_OFF = "FALSE",
    parameter integer PMA_REG_RX_ICTRL_EQ = 2,
    parameter PMA_REG_EQ_DC_CALIB_EN = "FALSE",
    parameter integer PMA_CTLE_CTRL_REG_I = 0,
    parameter PMA_CTLE_REG_FORCE_SEL_I = "FALSE",
    parameter PMA_CTLE_REG_HOLD_I = "FALSE",
    parameter integer PMA_CTLE_REG_INIT_DAC_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_INIT_DAC_I_3_2 = 0,
    parameter PMA_CTLE_REG_POLARITY_I = "FALSE",
    parameter integer PMA_CTLE_REG_SHIFTER_GAIN_I = 4,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_9_2 = 1,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_11_10 = 0,
    parameter PMA_REG_RX_RES_TRIM_EN = "FALSE",
    parameter integer PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION = 1,
    parameter integer PMA_REG_ALG_RX_TERM_VCM_SELECTION = 3,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0 = 0,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8 = 0,
    parameter PMA_REG_ALG_LOW_SPEED_MODE_ENABLE = "FALSE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER = "TRUE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION = "FALSE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_EYE_DFETAP1_PLORITY = "FALSE",
    parameter PMA_REG_CDR_SEL = "FALSE",
    parameter PMA_REG_EYE_DET_EN = "FALSE",
    parameter integer PMA_REG_PI_BIAS_CURRENT = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_6_0 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_14_7 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_21_15 = 0,
    parameter integer PMA_REG_ALG_EYE_PATH_SEL = 0,
    parameter integer PMA_REG_ALG_CTLE_TEST_SEL = 0,
    parameter PMA_REG_RX_SLIP_SEL_4 = "FALSE",
    parameter PMA_REG_ALG_RX_T1_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_CDRX_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_VP_T1_SW_PLORITY = "FALSE",
    parameter PMA_REG_ALG_RX_VP_PLORITY = "TRUE",
    parameter PMA_REG_ALG_RX_GAIN_CTRL_SUMMER = "FALSE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_T1_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_VP_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_EYE_EN = "TRUE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE = "FALSE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_REG = "FALSE",
    parameter PMA_REG_RX_PGA_OFF = "FALSE",
    parameter integer PMA_REG_ALG_CDR_XWEIGHT_I = 4,
    parameter integer PMA_REG_ALG_CDR_YWEIGHT_I = 4,
    parameter PMA_REG_ALG_CTLE_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_CTLE_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_CTLE_INITDAC_6 = 0,
    parameter PMA_REG_ALG_CTLE_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_2_0 = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_4_3 = 2,
    parameter PMA_REG_ALG_CTLEOFS_FLIPDIR_I = "TRUE",
    parameter PMA_REG_ALG_CTLEOFS_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_3_0 = 0,
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_6_4 = 4,
    parameter PMA_REG_ALG_CTLEOFS_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_SHIFT_I = 4,
    parameter PMA_REG_ALG_DFE_CTLE_PWD = "FALSE",
    parameter PMA_REG_ALG_H1_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H1_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_H1_INITDAC_6 = 0,
    parameter PMA_REG_ALG_H1_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_SHIFT_I = 4,
    parameter PMA_REG_ALG_H2_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H2_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H2_INITDAC_5_1 = 0,
    parameter PMA_REG_ALG_H2_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_SHIFT_I_1_0 = 0,
    parameter integer PMA_REG_ALG_H2_SHIFT_I_2 = 1,
    parameter PMA_REG_ALG_H3_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H3_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_INITDAC_4_0 = 0,
    parameter integer PMA_REG_ALG_H3_INITDAC_5 = 1,
    parameter PMA_REG_ALG_H3_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_SHIFT_I = 4,
    parameter PMA_REG_ALG_H4_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H4_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H4_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_H4_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_SHIFT_I = 4,
    parameter PMA_REG_ALG_H5_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H5_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_INITDAC = 16,
    parameter PMA_REG_ALG_H5_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_SHIFT_I = 4,
    parameter PMA_REG_ALG_H6_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H6_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_H6_INITDAC_4_3 = 2,
    parameter PMA_REG_ALG_H6_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_HCTLE_OFS_1_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OFS_3_2 = 2,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_6 = 1,
    parameter PMA_REG_ALG_HCTLE_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQH_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQH_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_REG_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_LEQL_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQL_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQL_REG_PRESELECT_I = 7,
    parameter integer PMA_REG_ALG_LEQL_REG_SHIFT_I = 4,
    parameter PMA_REG_ALG_NEXTBIT_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_6_0 = 127,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_14_7 = 255,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_19_15 = 31,
    parameter integer PMA_REG_ALG_SOFS_DACWIN_I = 1,
    parameter PMA_REG_ALG_SOFS_FLIP_DIR_I = "TRUE",
    parameter PMA_REG_ALG_SOFS_FORCE_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_5_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_6 = 1,
    parameter integer PMA_REG_ALG_SOFS_FORCENUM_I = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_6_3 = 8,
    parameter integer PMA_REG_ALG_SOFS_SHIFT_I = 1,
    parameter PMA_REG_ALG_SOFS_SKIP_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0 = 254,
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8 = 15,
    parameter PMA_REG_ALG_ST_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_ST_FORCEN = "FALSE",
    parameter PMA_REG_ALG_ST_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_ST_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_ST_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_ST_RECALEN = "FALSE",
    parameter integer PMA_REG_ALG_ST_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_ST_STARTCNT_7_0 = 0,
    parameter integer PMA_REG_ALG_ST_STARTCNT_15_8 = 128,
    parameter integer PMA_REG_ALG_ST_STARTCNT_19_16 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_3_0 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_11_4 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_17_12 = 2,
    parameter integer PMA_REG_ALG_ST_TOPTAP_1_0 = 3,
    parameter integer PMA_REG_ALG_ST_TOPTAP_3_2 = 3,
    parameter integer PMA_REG_ALG_SWCLK_DIV = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_3_0 = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_4 = 1,
    parameter integer PMA_REG_ALG_TAPA_NUM = 7,
    parameter integer PMA_REG_ALG_TAPB_DAC_0 = 0,
    parameter integer PMA_REG_ALG_TAPB_DAC_4_1 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_3_0 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_5_4 = 0,
    parameter integer PMA_REG_ALG_TAPC_DAC = 16,
    parameter integer PMA_REG_ALG_TAPC_NUM_0 = 1,
    parameter integer PMA_REG_ALG_TAPC_NUM_5_1 = 4,
    parameter integer PMA_REG_ALG_TAPD_DAC_2_0 = 0,
    parameter integer PMA_REG_ALG_TAPD_DAC_4_3 = 2,
    parameter integer PMA_REG_ALG_TAPD_NUM = 10,
    parameter PMA_REG_ALG_VP_FLIPDIR_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_GRN_SHIFT_I = 5,
    parameter PMA_REG_ALG_VP_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_IDEAL_2_0 = 0,
    parameter integer PMA_REG_ALG_VP_IDEAL_6_3 = 10,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_3_0 = 0,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_6_4 = 0,
    parameter PMA_REG_ALG_VP_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_VP_RED_SHIFT_I = 5,
    parameter integer PMA_REG_ALG_VPOFS_SEL_0 = 0,
    parameter integer PMA_REG_ALG_VPOFS_SEL_2_1 = 1,
    parameter integer PMA_REG_ALG_H1_UPBOUND_5_0 = 55,
    parameter integer PMA_REG_ALG_H1_UPBOUND_6 = 1,
    parameter PMA_REG_ALG_CTLEOFS_PWDN = "FALSE",
    parameter PMA_REG_ALG_LEQH_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_AGC_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_AGC_INITDAC = 10,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_1_0 = 3,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_3_2 = 0,
    parameter PMA_REG_ALG_AGC_OVERWREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_PWD = "FALSE",
    parameter integer PMA_REG_ALG_AGC_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_0 = 1,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_3_1 = 7,
    parameter integer PMA_REG_ALG_AGC_WAITSEL = 11,
    parameter PMA_REG_PI_CTRL_SEL_RX = "FALSE",
    parameter integer PMA_REG_PI_CTRL_RX_4_0 = 0,
    parameter integer PMA_REG_PI_CTRL_RX_7_5 = 0,
    parameter PMA_CFG_RX_LANE_POWERUP = "ON",
    parameter PMA_CFG_RX_PMA_RSTN = "TRUE",
    parameter PMA_INT_PMA_RX_MASK_0 = "FALSE",
    parameter PMA_INT_PMA_RX_CLR_0 = "FALSE",
    parameter PMA_CFG_CTLE_ADP_RSTN = "TRUE",
    parameter PMA_CFG_RX_CDR_RSTN = "TRUE",
    parameter PMA_CFG_RX_CLKPATH_RSTN = "TRUE",
    parameter PMA_CFG_RX_DFE_RSTN = "TRUE",
    parameter PMA_CFG_RX_LEQ_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIDING_RSTN = "TRUE",
    parameter PMA_CFG_RX_EYE_RSTN = "TRUE",
    parameter PMA_CFG_RX_CTLE_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLICER_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIP_RSTN = "TRUE",
    parameter integer PMA_REG_TX_BEACON_TIMER_SEL = 0,
    parameter PMA_REG_TX_BIT_CONV = "FALSE",
    parameter integer PMA_REG_TX_RES_CAL = 50,
    parameter integer PMA_REG_TX_UDP_DATA_20 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_26_21 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_34_27 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_39_25 = 0,
    parameter integer PMA_REG_TX_BUSWIDTH_EN = 0,
    parameter PMA_REG_TX_PD_POST = "OFF",
    parameter PMA_REG_TX_PD_POST_OW = "FALSE",
    parameter PMA_REG_TX_BUSWIDTH = "20BIT",
    parameter integer PMA_REG_EI_PCLK_DELAY_SEL = 0,
    parameter integer PMA_REG_TX_AMP_DAC0 = 25,
    parameter integer PMA_REG_TX_AMP_DAC1 = 19,
    parameter integer PMA_REG_TX_AMP_DAC2 = 14,
    parameter integer PMA_REG_TX_AMP_DAC3 = 9,
    parameter PMA_REG_TX_RXDET_THRESHOLD = "84MV",
    parameter PMA_REG_TX_BEACON_OSC_CTRL = "FALSE",
    parameter integer PMA_REG_TX_PRBS_GEN_WIDTH_SEL = 0,
    parameter PMA_REG_TX_TX2RX_SLPBACK_EN = "FALSE",
    parameter PMA_REG_TX_PCLK_EDGE_SEL = "FALSE",
    parameter PMA_REG_TX_PRBS_GEN_EN = "FALSE",
    parameter PMA_REG_TX_PRBS_SEL = "PRBS7",
    parameter integer PMA_REG_TX_UDP_DATA_7_TO_0 = 5,
    parameter integer PMA_REG_TX_UDP_DATA_15_TO_8 = 235,
    parameter integer PMA_REG_TX_UDP_DATA_19_TO_16 = 3,
    parameter integer PMA_REG_TX_FIFO_WP_CTRL = 4,
    parameter PMA_REG_TX_FIFO_EN = "FALSE",
    parameter integer PMA_REG_TX_DATA_MUX_SEL = 0,
    parameter PMA_REG_TX_ERR_INSERT = "FALSE",
    parameter PMA_REG_TX_SATA_EN = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON_OW = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON = "TRUE",
    parameter integer PMA_REG_TX_CFG_POST1 = 0,
    parameter integer PMA_REG_TX_CFG_POST2 = 0,
    parameter integer PMA_REG_TX_OOB_DELAY_SEL = 0,
    parameter PMA_REG_TX_POLARITY = "NORMAL",
    parameter PMA_REG_TX_LS_MODE_EN = "FALSE",
    parameter PMA_REG_RX_JTAG_OE = "TRUE",
    parameter integer PMA_REG_RX_ACJTAG_VHYSTSEL = 0,
    parameter PMA_REG_TX_RES_CAL_EN = "FALSE",
    parameter integer PMA_REG_RX_TERM_MODE_CTRL = 5,
    parameter PMA_REG_PLPBK_TXPCLK_EN = "FALSE",
    parameter integer PMA_REG_CLK_SEL_STROBE_TXPCLK = 2,
    parameter integer PMA_REG_TX_PH_SEL_0 = 1,
    parameter integer PMA_REG_TX_PH_SEL_6_1 = 0,
    parameter integer PMA_REG_TX_CFG_PRE = 0,
    parameter integer PMA_REG_TX_CFG_MAIN = 0,
    parameter integer PMA_REG_CFG_POST = 0,
    parameter PMA_REG_PD_MAIN = "TRUE",
    parameter PMA_REG_PD_PRE = "TRUE",
    parameter integer PMA_REG_TX_RXDET_TIMER_SEL = 87,
    parameter PMA_REG_TX_PI_CUR_BUF = "10GHz",
    parameter PMA_REG_TX_MOD_STAND_BY_EN = "FALSE",
    parameter PMA_REG_STATE_STAND_BY_SEL = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_POLAR_CTRL = "FALSE",
    parameter PMA_REG_TX_FREERUN_PD = "TRUE",
    parameter PMA_REG_TX_CHANGE_ON_SEL = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_CTRL = "FALSE",
    parameter integer PMA_REG_TX_FREERUN_RATE_0 = 0,
    parameter integer PMA_REG_TX_FREERUN_RATE_1 = 0,
    parameter PMA_REG_TX_FREERUN_RATE_OW = "FALSE",
    parameter PMA_REG_TX_RST_SYNC_CLK_SEL = "TRUE",
    parameter integer PMA_REG_TX_PI_CTRL_SEL = 0,
    parameter integer PMA_REG_TX_PI_CTRL = 0,
    parameter PMA_LANE_POWERUP = "TRUE",
    parameter PMA_POR_N = "TRUE",
    parameter PMA_TX_LANE_POWERUP = "TRUE",
    parameter PMA_TX_PMA_RSTN = "TRUE",
    parameter PMA_LPLL_POWERUP = "TRUE",
    parameter PMA_LPLL_RSTN = "TRUE",
    parameter PMA_LPLL_LOCKDET_RSTN = "TRUE",
    parameter integer PMA_REG_LPLL_PFDDELAY_SEL = 1,
    parameter PMA_REG_LPLL_PFDDELAY_EN = "TRUE",
    parameter integer PMA_REG_LPLL_VCTRL_SET = 0,
    parameter PMA_LPLL_CHARGE_PUMP_CTRL = "type",
    parameter PMA_LPLL_REFDIV = "DIV1",
    parameter integer PMA_LPLL_FBDIV = 38,
    parameter integer PMA_LPLL_LPF_RES = 1,
    parameter integer PMA_LPLL_REFLOSS_READY = 0,
    parameter integer PMA_LPLL_LOCKED_PFDDELAY = 0,
    parameter integer PMA_LPLL_MCLK_SEL = 0,
    parameter integer PMA_LPLL_TEST_SEL = 0,
    parameter PMA_LPLL_TEST_SIG_HALF_EN = "TRUE",
    parameter PMA_LPLL_TEST_V_EN = "FALSE",
    parameter PMA_LPLL_MCLK_EN = "TRUE",
    parameter integer PMA_LPLL_MCLK_DET_CTL = 16,
    parameter integer PMA_LPLL_LOCKDET_REFCT = 3,
    parameter integer PMA_LPLL_LOCKDET_FBCT = 3,
    parameter integer PMA_LPLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_LPLL_LOCKDET_ITER = 1,
    parameter integer PMA_LPLL_UNLOCKDET_ITER = 2,
    parameter integer PMA_LPLL_LOCKDET_EN_OW = 0,
    parameter integer PMA_LPLL_LOCKDET_EN = 0,
    parameter integer PMA_LPLL_LOCKDET_MODE = 0,
    parameter integer PMA_LPLL_LOCKDET_OW = 0,
    parameter integer PMA_LPLL_LOCKDETED = 0,
    parameter integer PMA_LPLL_UNLOCKDET_OW = 0,
    parameter integer PMA_LPLL_UNLOCKDETED = 0,
    parameter integer PMA_LPLL_LOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_UNLOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_LOCKDET_REPEAT = 0,
    parameter integer PMA_LPLL_NOFBCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_NOREFCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_READY_OR_LOCK = 0,
    parameter integer PMA_LPLL_READY = 0,
    parameter integer PMA_LPLL_READY_OW = 0,
    parameter PMA_REG_TXCLK_SEL = "HPLL",
    parameter PMA_REG_RXCLK_SEL = "HPLL",
    parameter integer PMA_REG_TEST_BUF = 0,
    parameter PMA_REG_RX_DEF_SEL0 = "18.75uA",
    parameter PMA_REG_RX_DEF_SEL1 = "18.75uA",
    parameter PMA_REG_TX_DIV_SEL = "25uA",
    parameter PMA_REG_LPLL_AMP_SEL = "25uA",
    parameter PMA_REG_LPLL_VCO_SEL = "25uA",
    parameter PMA_REG_LPLL_CHARGE_PUMP_SEL = "25uA",
    parameter PMA_REG_RX_EQ0_SEL = "56.25uA",
    parameter PMA_REG_RX_EQ1_SEL = "56.25uA",
    parameter PMA_REG_RX_PGA_SEL = "56.25uA",
    parameter integer PMA_REG_CHL_TEST = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_7_0 = 255,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_15_8 = 247,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_18_16 = 7,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_21_19 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_29_22 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_37_30 = 1,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_4_0 = 31,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_8_5 = 15,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_12_9 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_17_13 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0
) (
    output P_CFG_READY,
    output [7:0] P_CFG_RDATA,
    output P_CFG_INT,
    output [24:0] LANE_COUT_BUS_FORWARD,
    output [1:0] LANE_COUT_BUS_BACKWARD,
    output P_RX_PRBS_ERROR,
    output P_PCS_RX_MCB_STATUS,
    output P_PCS_LSM_SYNCED,
    output [87:0] P_RDATA,
    output P_RXDVLD,
    output P_RXDVLD_H,
    output [5:0] P_RXSTATUS,
    output [2:0] P_EM_ERROR_CNT,
    output P_LPLL_READY,
    output P_RX_SIGDET_STATUS,
    output P_RX_SATA_COMINIT,
    output P_RX_SATA_COMWAKE,
    output P_RX_LS_DATA,
    output P_RX_READY,
    output [19:0] P_TEST_STATUS,
    output P_TX_RXDET_STATUS,
    output P_RCLK2FABRIC,
    output P_TCLK2FABRIC,
    output P_CA_ALIGN_RX,
    output P_CA_ALIGN_TX,
    output P_TX_SDN,
    output P_TX_SDP,
    input P_RX_CLK_FR_CORE,
    input P_RCLK2_FR_CORE,
    input P_TX_CLK_FR_CORE,
    input P_TCLK2_FR_CORE,
    input P_PCS_RX_RST,
    input P_PCS_TX_RST,
    input P_EXT_BRIDGE_PCS_RST,
    input P_CFG_RST,
    input P_CFG_CLK,
    input P_CFG_PSEL,
    input P_CFG_ENABLE,
    input P_CFG_WRITE,
    input [11:0] P_CFG_ADDR,
    input [7:0] P_CFG_WDATA,
    input [24:0] LANE_CIN_BUS_FORWARD,
    input [1:0] LANE_CIN_BUS_BACKWARD,
    input [87:0] P_TDATA,
    input P_PCIE_EI_H,
    input P_PCIE_EI_L,
    input [15:0] P_TX_DEEMP,
    input [1:0] P_TX_DEEMP_POST_SEL,
    input P_BLK_ALIGN_CTRL,
    input P_TX_ENC_TYPE,
    input P_RX_DEC_TYPE,
    input P_PCS_BIT_SLIP,
    input P_PCS_WORD_ALIGN_EN,
    input P_RX_POLARITY_INVERT,
    input P_PCS_MCB_EXT_EN,
    input P_PCS_NEAREND_LOOP,
    input P_PCS_FAREND_LOOP,
    input P_PMA_NEAREND_PLOOP,
    input P_PMA_NEAREND_SLOOP,
    input P_PMA_FAREND_PLOOP,
    input P_PCS_PRBS_EN,
    input P_LANE_POWERDOWN,
    input P_LANE_RST,
    input P_RX_LANE_POWERDOWN,
    input P_RX_PMA_RST,
    input P_RX_CDR_RST,
    input P_RX_CLKPATH_RST,
    input P_RX_DFE_RST,
    input P_RX_LEQ_RST,
    input P_RX_SLIDING_RST,
    input P_RX_DFE_EN,
    input P_RX_T1_EN,
    input P_RX_CDRX_EN,
    input P_RX_T1_DFE_EN,
    input P_RX_T2_DFE_EN,
    input P_RX_T3_DFE_EN,
    input P_RX_T4_DFE_EN,
    input P_RX_T5_DFE_EN,
    input P_RX_T6_DFE_EN,
    input P_RX_SLIDING_EN,
    input P_RX_EYE_RST,
    input P_RX_EYE_EN,
    input [7:0] P_RX_EYE_TAP,
    input [7:0] P_RX_PIC_EYE,
    input [7:0] P_RX_PIC_FASTLOCK,
    input P_RX_PIC_FASTLOCK_STROBE,
    input P_EM_RD_TRIGGER,
    input [1:0] P_EM_MODE_CTRL,
    input P_RX_CTLE_DCCAL_RST,
    input P_RX_SLICER_DCCAL_RST,
    input P_RX_SLICER_DCCAL_EN,
    input P_RX_CTLE_DCCAL_EN,
    input P_RX_SLIP_RST,
    input P_RX_SLIP_EN,
    input P_LPLL_POWERDOWN,
    input P_LPLL_RST,
    input P_LPLL_LOCKDET_RST,
    input P_TX_LS_DATA,
    input P_TX_BEACON_EN,
    input P_TX_SWING,
    input P_TX_RXDET_REQ,
    input [1:0] P_TX_RATE,
    input [2:0] P_TX_BUSWIDTH,
    input [2:0] P_TX_FREERUN_BUSWIDTH,
    input [2:0] P_TX_MARGIN,
    input P_TX_PMA_RST,
    input P_TX_LANE_POWERDOWN,
    input P_TX_PIC_EN,
    input [1:0] P_RX_RATE,
    input [2:0] P_RX_BUSWIDTH,
    input P_RX_HIGHZ,
    input [7:0] P_CIM_CLK_ALIGNER_RX,
    input [7:0] P_CIM_CLK_ALIGNER_TX,
    input P_ALIGN_MODE_VALID_RX,
    input [1:0] P_ALIGN_MODE_RX,
    input P_ALIGN_MODE_VALID_TX,
    input [2:0] P_ALIGN_MODE_TX,
    input PMA_HPLL_CK0,
    input PMA_HPLL_CK90,
    input PMA_HPLL_CK180,
    input PMA_HPLL_CK270,
    input PMA_HPLL_READY_IN,
    input PMA_HPLL_REFCLK_IN,
    input PMA_TX_SYNC_HPLL_IN,
    input P_LPLL_REFCLK_IN,
    input P_TX_RATE_CHANGE_ON_0,
    input P_TX_RATE_CHANGE_ON_1,
    input P_TX_SYNC,
    input P_RX_SDN,
    input P_RX_SDP,
    output P_TEST_SO0,
    output P_TEST_SO1,
    output P_TEST_SO2,
    output P_TEST_SO3,
    output P_TEST_SO4,
    output [1:0] P_FOR_PMA_TEST_SO,
    input P_TEST_SE_N,
    input P_TEST_MODE_N,
    input P_TEST_RSTN,
    input P_TEST_SI0,
    input P_TEST_SI1,
    input P_TEST_SI2,
    input P_TEST_SI3,
    input P_TEST_SI4,
    input P_FOR_PMA_TEST_MODE_N,
    input [1:0] P_FOR_PMA_TEST_SE_N,
    input [1:0] P_FOR_PMA_TEST_CLK,
    input [1:0] P_FOR_PMA_TEST_RSTN,
    input [1:0] P_FOR_PMA_TEST_SI
)  ;
endmodule


module GTP_HSSTHP_LANE_E1
#(
    parameter PCS_DYN_DLY_SEL_RX = "FALSE",
    parameter PCS_PMA_RCLK_POLINV = "PMA_RCLK",
    parameter PCS_PCS_RCLK_SEL = "RCLK",
    parameter PCS_GEAR_RCLK_SEL = "RCLK",
    parameter PCS_RCLK2FABRIC_SEL = "HARD_1",
    parameter PCS_SCAN_INTERVAL_RX = "4_CLOCKS",
    parameter PCS_BRIDGE_RCLK_SEL = "RCLK",
    parameter PCS_RCLK_POLINV = "RCLK",
    parameter PCS_TO_FABRIC_CLK_SEL = "PMA_RCLK",
    parameter PCS_CLK2ALIGNER_SEL = "TO_FABRIC_CLK",
    parameter PCS_TO_FABRIC_CLK_DIV_EN = "FALSE",
    parameter PCS_AUTO_NEAR_LOOP_EN = "FALSE",
    parameter PCS_PCS_RCLK_EN = "FALSE",
    parameter PCS_BRIDGE_PCS_RCLK_EN_SEL = "HARD_1",
    parameter PCS_BRIDGE_RCLK_EN_SEL = "HARD_0",
    parameter PCS_GEAR_RCLK_EN_SEL = "HARD_0",
    parameter PCS_NEGEDGE_EN_RX = "FALSE",
    parameter PCS_PCS_RX_RSTN = "FALSE",
    parameter PCS_BRIDGE_PCS_RSTN = "FALSE",
    parameter PCS_TO_FABRIC_RST_EN = "FALSE",
    parameter PCS_BYPASS_GEAR_RRSTN = "FALSE",
    parameter PCS_BYPASS_BRIDGE_RRSTN = "FALSE",
    parameter PCS_ALIGNER_EN_RX = "FALSE",
    parameter PCS_RX_SLAVE = "MASTER",
    parameter integer PCS_RX_CA = 0,
    parameter integer PCS_SUM_THRESHOLD_RX = 0,
    parameter integer PCS_AVG_CYCLES_RX = 0,
    parameter PCS_REG_PMA_RX2TX_PLOOP_EN = "FALSE",
    parameter PCS_REG_PMA_RX2TX_PLOOP_FIFOEN = "FALSE",
    parameter integer PCS_STEP_SIZE_RX = 0,
    parameter integer PCS_REV_CNT_LIMIT_RX = 0,
    parameter integer PCS_FILTER_CNT_SIZE_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_3_0 = 0,
    parameter integer PCS_DLY_REC_SIZE_RX = 0,
    parameter integer PCS_ALIGN_THRD_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_4 = 0,
    parameter PCS_CFG_DEC_TYPE_EN = "FALSE",
    parameter PCS_RXBRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_GE_AUTO_EN = "FALSE",
    parameter PCS_RXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_RXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_IFG_EN = "FALSE",
    parameter PCS_FLP_FULL_CHK_EN = "FALSE",
    parameter PCS_FLP_EMPTY_CHK_EN = "FALSE",
    parameter PCS_RX_POLARITY_INV = "DELAY",
    parameter PCS_FARLP_PWR_REDUCTION = "FALSE",
    parameter PCS_RXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_WDALIGN_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXDEC_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXTEST_PWR_REDUCTION = "NORMAL",
    parameter integer PCS_WA_SOS_DET_TOL = 0,
    parameter integer PCS_WA_SE_DET_TOL = 0,
    parameter PCS_RX_SAMPLE_UNION = "FALSE",
    parameter PCS_NEAR_LOOP = "FALSE",
    parameter PCS_BYPASS_WORD_ALIGN = "FALSE",
    parameter PCS_BYPASS_DENC = "FALSE",
    parameter PCS_RX_ERRCNT_CLR = "FALSE",
    parameter PCS_RX_CODE_MODE = "DUAL_8B10B",
    parameter PCS_RX_BYPASS_GEAR = "FALSE",
    parameter PCS_ERRDETECT_SILENCE = "FALSE",
    parameter PCS_RX_DATA_MODE = "8BIT",
    parameter PCS_CA_DYN_CLY_EN_RX = "FALSE",
    parameter PCS_CFG_APATTERN_STATUS_DELAY = "DELAY_ONE_CYCLE",
    parameter PCS_RX_PRBS_MODE = "DISABLE",
    parameter PCS_ALIGN_MODE = "1GB",
    parameter PCS_COMMA_DET_MODE = "PATTERN_DETECT",
    parameter integer PCS_RAPID_VMIN_1 = 0,
    parameter integer PCS_RAPID_VMIN_2 = 0,
    parameter PCS_RXBU_WIDER_EN = "40/20BIT",
    parameter integer PCS_RAPID_IMAX = 0,
    parameter PCS_RX_SPLIT = "SPLIT_22BIT_11BIT",
    parameter integer PCS_RXBRG_END_PACKET_9_8 = 0,
    parameter integer PCS_RXBRG_END_PACKET_7_0 = 0,
    parameter integer PCS_CTC_MAX_DEL = 0,
    parameter integer PCS_COMMA_REG0_9_8 = 0,
    parameter integer PCS_COMMA_REG1_9_8 = 0,
    parameter integer PCS_COMMA_MASK_9_8 = 0,
    parameter integer PCS_COMMA_REG0_7_0 = 0,
    parameter integer PCS_COMMA_REG1_7_0 = 0,
    parameter integer PCS_COMMA_MASK_7_0 = 0,
    parameter integer PCS_FLP_WRADDR_START = 0,
    parameter integer PCS_FLP_RDADDR_START = 0,
    parameter PCS_CFG_RX_BRIDGE_CLK_POLINV = "FALSE",
    parameter PCS_CTC_MODE_RD_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AFULL = 0,
    parameter PCS_FAST_LOCK_GEAR_EN = "FALSE",
    parameter PCS_CTC_MODE_WR_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AEMPTY = 0,
    parameter PCS_CTC_MODE = "ONE_BYTE",
    parameter PCS_RXBRIDGE_MODE = "BYPASS",
    parameter integer PCS_CTC_ADD_MAX = 0,
    parameter PCS_CFG_PHDET_EN_RX = "FALSE",
    parameter integer PCS_WA_SDS_DET_TOL = 0,
    parameter PCS_CEB_MODE = "10GB",
    parameter PCS_APATTERN_MODE = "ONE_BYTE",
    parameter PCS_A_REG0_8 = "FALSE",
    parameter integer PCS_RXBRG_WADDR_START = 0,
    parameter PCS_A_REG1_8 = "FALSE",
    parameter integer PCS_RXBRG_RADDR_START = 0,
    parameter integer PCS_A_REG0_7_0 = 0,
    parameter integer PCS_A_REG1_7_0 = 0,
    parameter integer PCS_CEB_RAPIDLS_MMAX = 0,
    parameter integer PCS_CEB_DETECT_TIME = 0,
    parameter integer PCS_WL_FIFO_RD = 0,
    parameter integer PCS_SKIP_REG0_9_8 = 0,
    parameter integer PCS_SKIP_REG0_7_0 = 0,
    parameter integer PCS_CFG_CONTI_SKP_SET = 0,
    parameter PCS_CFG_RX_BASE_ADV_MODE = "BASE_MODE",
    parameter integer PCS_SKIP_REG1_9_8 = 0,
    parameter integer PCS_SKIP_REG2_9_8 = 0,
    parameter integer PCS_SKIP_REG3_9_8 = 0,
    parameter integer PCS_SKIP_REG1_7_0 = 0,
    parameter integer PCS_SKIP_REG2_7_0 = 0,
    parameter integer PCS_SKIP_REG3_7_0 = 0,
    parameter integer PCS_CFG_PRBS_ERR_O_SEL = 0,
    parameter integer PCS_CFG_PD_DELAY_RX = 0,
    parameter integer PCS_WR_START_GAP = 0,
    parameter integer PCS_MIN_IFG = 0,
    parameter PCS_INT_RX_MASK_0 = "FALSE",
    parameter PCS_INT_RX_MASK_1 = "FALSE",
    parameter PCS_INT_RX_MASK_2 = "FALSE",
    parameter PCS_INT_RX_MASK_3 = "FALSE",
    parameter PCS_INT_RX_MASK_4 = "FALSE",
    parameter PCS_INT_RX_MASK_5 = "FALSE",
    parameter PCS_INT_RX_CLR_5 = "FALSE",
    parameter PCS_INT_RX_CLR_4 = "FALSE",
    parameter PCS_INT_RX_CLR_3 = "FALSE",
    parameter PCS_INT_RX_CLR_2 = "FALSE",
    parameter PCS_INT_RX_CLR_1 = "FALSE",
    parameter PCS_INT_RX_CLR_0 = "FALSE",
    parameter PCS_EM_CNT_RD_EN = "FALSE",
    parameter PCS_EM_CTRL_SEL = "SIGNAL_CTRL",
    parameter PCS_EM_MODE_CTRL = "HOLD",
    parameter PCS_EM_RD_CONDITION = "TRIGGER",
    parameter integer PCS_EM_SP_PATTERN_7_0 = 0,
    parameter integer PCS_EM_SP_PATTERN_15_8 = 0,
    parameter integer PCS_EM_SP_PATTERN_23_16 = 0,
    parameter integer PCS_EM_SP_PATTERN_31_24 = 0,
    parameter integer PCS_EM_SP_PATTERN_39_32 = 0,
    parameter integer PCS_EM_SP_PATTERN_47_40 = 0,
    parameter integer PCS_EM_SP_PATTERN_55_48 = 0,
    parameter integer PCS_EM_SP_PATTERN_63_56 = 0,
    parameter integer PCS_EM_SP_PATTERN_71_64 = 0,
    parameter integer PCS_EM_SP_PATTERN_79_72 = 0,
    parameter integer PCS_EM_PMA_MASK_7_0 = 0,
    parameter integer PCS_EM_PMA_MASK_15_8 = 0,
    parameter integer PCS_EM_PMA_MASK_23_16 = 0,
    parameter integer PCS_EM_PMA_MASK_31_24 = 0,
    parameter integer PCS_EM_PMA_MASK_39_32 = 0,
    parameter integer PCS_EM_PMA_MASK_47_40 = 0,
    parameter integer PCS_EM_PMA_MASK_55_48 = 0,
    parameter integer PCS_EM_PMA_MASK_63_56 = 0,
    parameter integer PCS_EM_PMA_MASK_71_64 = 0,
    parameter integer PCS_EM_PMA_MASK_79_72 = 0,
    parameter integer PCS_EM_EYED_MASK_7_0 = 0,
    parameter integer PCS_EM_EYED_MASK_15_8 = 0,
    parameter integer PCS_EM_EYED_MASK_23_16 = 0,
    parameter integer PCS_EM_EYED_MASK_31_24 = 0,
    parameter integer PCS_EM_EYED_MASK_39_32 = 0,
    parameter integer PCS_EM_EYED_MASK_47_40 = 0,
    parameter integer PCS_EM_EYED_MASK_55_48 = 0,
    parameter integer PCS_EM_EYED_MASK_63_56 = 0,
    parameter integer PCS_EM_EYED_MASK_71_64 = 0,
    parameter integer PCS_EM_EYED_MASK_79_72 = 0,
    parameter integer PCS_EM_PRESCALE = 0,
    parameter PCS_CFG_TEST_STATUS_SEL = "SEL_PMA_TEST_STATUS_INT",
    parameter integer PCS_CFG_DIFF_CNT_BND_RX = 0,
    parameter PCS_CFG_FLT_SEL_RX = "FALSE",
    parameter integer PCS_FILTER_BND_RX = 0,
    parameter PCS_TCLK2FABRIC_DIV_RST_M = "FALSE",
    parameter PCS_TX_PMA_TCLK_POLINV = "PMA_TCLK",
    parameter PCS_TX_TCLK_POLINV = "TCLK",
    parameter PCS_PCS_TCLK_SEL = "PMA_TCLK",
    parameter PCS_GEAR_TCLK_SEL = "PMA_TCLK",
    parameter PCS_TX_BRIDGE_TCLK_SEL = "TCLK",
    parameter PCS_TCLK2ALIGNER_SEL = "PMA_TCLK",
    parameter CA_DYN_DLY_EN_TX = "FALSE",
    parameter PCS_TX_PCS_CLK_EN_SEL = "HARDWIRED1",
    parameter PCS_TX_GEAR_CLK_EN_SEL = "HARDWIRED0",
    parameter PCS_TCLK2FABRIC_DIV_EN = "FALSE",
    parameter PCS_TCLK2FABRIC_SEL = "CLK2ALIGNER_N_DIV2",
    parameter integer DLY_ADJUST_SIZE_TX = 0,
    parameter PCS_TX_PCS_TX_RSTN = "FALSE",
    parameter PCS_TX_CA_RSTN = "FALSE",
    parameter PCS_TX_SLAVE = "MASTER",
    parameter integer PCS_TX_CA = 0,
    parameter integer PCS_CFG_PI_CLK_SEL = 0,
    parameter PCS_CFG_PI_CLK_EN_SEL = "CLK_EN_ALWAYS1",
    parameter integer PCS_CFG_PI_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_SUM_THRESHOLD_TX = 0,
    parameter integer PCS_CFG_AVG_CYCLES_TX = 0,
    parameter PCS_CFG_NEGEDGE_EN_TX = "FALSE",
    parameter integer PCS_CFG_ALIGN_THRD_TX = 0,
    parameter integer PCS_CFG_SCAN_INTERVAL_TX = 0,
    parameter integer PCS_CFG_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_REV_CNT_LIMIT_TX = 0,
    parameter integer PCS_CFG_FILTER_CNT_SIZE_TX = 0,
    parameter integer PCS_CFG_PI_DEFAULT_TX = 0,
    parameter PCS_CFG_PHDET_EN_TX = "FALSE",
    parameter PCS_PMA_TX2RX_PLOOP_EN = "FALSE",
    parameter PCS_PMA_TX2RX_SLOOP_EN = "FALSE",
    parameter PCS_CFG_DYN_DLY_SEL_TX = "FALSE",
    parameter integer PCS_CFG_DLY_REC_SIZE_TX = 0,
    parameter PCS_TX_DATA_WIDTH_MODE = "8BIT",
    parameter PCS_TX_BYPASS_BRIDGE_UINT = "FALSE",
    parameter PCS_TX_BYPASS_BRIDGE_FIFO = "FALSE",
    parameter PCS_TX_BYPASS_GEAR = "FALSE",
    parameter PCS_TX_BYPASS_ENC = "FALSE",
    parameter PCS_TX_BYPASS_BIT_SLIP = "FALSE",
    parameter PCS_TX_BRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_TXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXGEAR_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXENC_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBSLP_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_TXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_TX_ENCODER_MODE = "DUAL_8B10B",
    parameter PCS_TX_PRBS_MODE = "DISABLE",
    parameter PCS_TX_DRIVE_REG_MODE = "NO_CHANGE",
    parameter integer PCS_TX_BIT_SLIP_CYCLES = 0,
    parameter PCS_TX_BASE_ADV_MODE = "BASE",
    parameter PCS_TX_GEAR_SPLIT = "NO_SPILT",
    parameter PCS_RX_BRIDGE_CLK_POLINV = "N_CLK_INVERT",
    parameter PCS_PRBS_ERR_LPBK = "FALSE",
    parameter PCS_TX_INSERT_ER = "FALSE",
    parameter PCS_ENABLE_PRBS_GEN = "FALSE",
    parameter PCS_FAR_LOOP = "FALSE",
    parameter PCS_CFG_ENC_TYPE_EN = "FALSE",
    parameter integer PCS_TXBRG_WADDR_START = 0,
    parameter integer PCS_TXBRG_RADDR_START = 0,
    parameter PCS_CFG_TX_PIC_EN = "DISABLE",
    parameter PCS_CFG_PIC_DIRECT_INV = "FALSE",
    parameter PCS_CFG_PI_MOD_CLK_EN = "FALSE",
    parameter PCS_CFG_TX_MODULATOR_OW_EN = "FALSE",
    parameter PCS_CFG_TX_PI_SSC_MODE_EN = "FALSE",
    parameter PCS_CFG_TX_PI_OFFSET_MODE_EN = "FALSE",
    parameter integer PCS_CFG_TX_PI_SSC_MODE_SEL = 0,
    parameter PCS_CFG_TXDEEMPH_EN = "FALSE",
    parameter PCS_PI_STROBE_SEL = "FALSE",
    parameter PCS_CFG_TX_PIC_GREY_SEL = "FALSE",
    parameter PCS_CFG_PIC_RENEW_INV = "NORMAL",
    parameter integer PCS_CFG_NUM_PIC = 0,
    parameter PCS_CFG_TXPIC_OW_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_OW_VALUE_0_7 = 0,
    parameter PCS_INT_TX_MASK_0 = "FALSE",
    parameter PCS_INT_TX_MASK_1 = "FALSE",
    parameter PCS_INT_TX_MASK_2 = "FALSE",
    parameter PCS_TX_WPTR_SEL = "FALSE",
    parameter PCS_INT_TX_CLR_2 = "FALSE",
    parameter PCS_INT_TX_CLR_1 = "FALSE",
    parameter PCS_INT_TX_CLR_0 = "FALSE",
    parameter integer PCS_CFG_PD_DELAY_TX = 0,
    parameter integer PCS_CFG_DIFF_CNT_BND_TX = 0,
    parameter PCS_CFG_PD_CLK_FR_CORE_SEL = "FALSE",
    parameter PCS_CFG_FLT_SEL_TX = "FALSE",
    parameter integer PCS_FILTER_BND_TX = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_7_0 = 0,
    parameter PCS_CFG_TX_SSC_MODULATOR_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_SCALE2_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_SCALE_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_8_9 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_8 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_8_9 = 0,
    parameter PMA_REG_CHL_BIAS_POWER_SEL = "FALSE",
    parameter PMA_REG_CHL_BIAS_POWER = "FALSE",
    parameter PMA_REG_RX_BUSWIDTH = "40BIT",
    parameter PMA_REG_RX_RATE = "DIV4",
    parameter PMA_REG_RX_RATE_EN = "FALSE",
    parameter integer PMA_REG_RX_RES_TRIM = 55,
    parameter PMA_REG_RX_SIGDET_STATUS_EN = "FALSE",
    parameter integer PMA_REG_CDR_READY_THD_7_0 = 32,
    parameter integer PMA_REG_CDR_READY_THD_11_8 = 0,
    parameter PMA_REG_RX_BUSWIDTH_EN = "FALSE",
    parameter PMA_REG_RX_PCLK_EDGE_SEL = "POS_EDGE",
    parameter integer PMA_REG_RX_PIBUF_IC = 3,
    parameter integer PMA_REG_RX_DCC_IC_RX = 1,
    parameter integer PMA_REG_CDR_READY_CHECK_CTRL = 0,
    parameter PMA_REG_RX_ICTRL_TRX = "100PCT",
    parameter integer PMA_REG_PRBS_CHK_WIDTH_SEL = 1,
    parameter PMA_REG_RX_ICTRL_PIBUF = "100PCT",
    parameter PMA_REG_RX_ICTRL_PI = "100PCT",
    parameter PMA_REG_RX_ICTRL_DCC = "100PCT",
    parameter PMA_REG_TX_RATE = "DIV1",
    parameter PMA_REG_TX_RATE_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N = "TRUE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_EN = "FALSE",
    parameter PMA_REG_RX_DATA_POLARITY = "NORMAL",
    parameter PMA_REG_RX_ERR_INSERT = "FALSE",
    parameter PMA_REG_UDP_CHK_EN = "FALSE",
    parameter PMA_REG_PRBS_SEL = "PRBS7",
    parameter PMA_REG_PRBS_CHK_EN = "FALSE",
    parameter integer PMA_REG_LPLL_NFC_STIC_DIS_N = 0,
    parameter PMA_REG_BIST_CHK_PAT_SEL = "PRBS",
    parameter PMA_REG_LOAD_ERR_CNT = "FALSE",
    parameter PMA_REG_CHK_COUNTER_EN = "TRUE",
    parameter integer PMA_REG_CDR_PROP_GAN_SEL = 3,
    parameter integer PMA_REG_CDR_TUBO_PROP_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_GAIN_SEL = 2,
    parameter integer PMA_REG_CDR_TUBO_INT_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_4_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_9_5 = 28,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_2_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_9_3 = 16,
    parameter integer PMA_ANA_RX_REG_O_61_55 = 21,
    parameter integer PMA_ANA_RX_REG_O_69_62 = 0,
    parameter integer PMA_ANA_RX_REG_O_77_70 = 135,
    parameter integer PMA_ANA_RX_REG_O_85_78 = 1,
    parameter integer PMA_ANA_RX_REG_O_93_86 = 8,
    parameter integer PMA_ANA_RX_REG_O_100_94 = 64,
    parameter integer PMA_ANA_RX_REG_O_108_101 = 0,
    parameter integer PMA_ANA_RX_REG_O_111_109 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_4_0 = 3,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_5 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MAX = 11,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MIN = 15,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MAX = 35,
    parameter integer PMA_REG_COMWAKE_STATUS_CLEAR = 0,
    parameter integer PMA_REG_COMINIT_STATUS_CLEAR = 0,
    parameter PMA_REG_RX_SATA_COMINIT_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMINIT = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE = "FALSE",
    parameter PMA_REG_RX_DCC_DISABLE = "FALSE",
    parameter PMA_REG_RX_SLIP_SEL_EN = "FALSE",
    parameter integer PMA_REG_RX_SLIP_SEL_3_0 = 0,
    parameter PMA_REG_RX_SLIP_EN = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_STATUS_SEL = 5,
    parameter PMA_REG_RX_SIGDET_FSM_RST_N = "TRUE",
    parameter PMA_REG_RX_SIGDET_STATUS = "FALSE",
    parameter PMA_REG_RX_SIGDET_VTH = "36MV",
    parameter integer PMA_REG_RX_SIGDET_GRM = 0,
    parameter PMA_REG_RX_SIGDET_PULSE_EXT = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_CH2_SEL = 0,
    parameter integer PMA_REG_RX_SIGDET_CH2_CHK_WINDOW = 3,
    parameter PMA_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",
    parameter integer PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0 = 0,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3 = 0,
    parameter integer PMA_REG_RX_SIGDET_4OOB_DET_SEL = 7,
    parameter integer PMA_REG_RX_SIGDET_IC_I = 10,
    parameter integer PMA_REG_RX_EQ1_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ1_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ1_OFF = "FALSE",
    parameter integer PMA_REG_RX_EQ2_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ2_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ2_OFF = "FALSE",
    parameter integer PMA_REG_RX_ICTRL_EQ = 2,
    parameter PMA_REG_EQ_DC_CALIB_EN = "FALSE",
    parameter integer PMA_CTLE_CTRL_REG_I = 0,
    parameter PMA_CTLE_REG_FORCE_SEL_I = "FALSE",
    parameter PMA_CTLE_REG_HOLD_I = "FALSE",
    parameter integer PMA_CTLE_REG_INIT_DAC_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_INIT_DAC_I_3_2 = 0,
    parameter PMA_CTLE_REG_POLARITY_I = "FALSE",
    parameter integer PMA_CTLE_REG_SHIFTER_GAIN_I = 4,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_9_2 = 1,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_11_10 = 0,
    parameter PMA_REG_RX_RES_TRIM_EN = "FALSE",
    parameter integer PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION = 1,
    parameter integer PMA_REG_ALG_RX_TERM_VCM_SELECTION = 3,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0 = 0,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8 = 0,
    parameter PMA_REG_ALG_LOW_SPEED_MODE_ENABLE = "FALSE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER = "TRUE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION = "FALSE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_EYE_DFETAP1_PLORITY = "FALSE",
    parameter PMA_REG_CDR_SEL = "FALSE",
    parameter PMA_REG_EYE_DET_EN = "FALSE",
    parameter integer PMA_REG_PI_BIAS_CURRENT = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_6_0 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_14_7 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_21_15 = 0,
    parameter integer PMA_REG_ALG_EYE_PATH_SEL = 0,
    parameter integer PMA_REG_ALG_CTLE_TEST_SEL = 0,
    parameter PMA_REG_RX_SLIP_SEL_4 = "FALSE",
    parameter PMA_REG_ALG_RX_T1_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_CDRX_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_VP_T1_SW_PLORITY = "FALSE",
    parameter PMA_REG_ALG_RX_VP_PLORITY = "TRUE",
    parameter PMA_REG_ALG_RX_GAIN_CTRL_SUMMER = "FALSE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_T1_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_VP_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_EYE_EN = "TRUE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE = "FALSE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_REG = "FALSE",
    parameter PMA_REG_RX_PGA_OFF = "FALSE",
    parameter integer PMA_REG_ALG_CDR_XWEIGHT_I = 4,
    parameter integer PMA_REG_ALG_CDR_YWEIGHT_I = 4,
    parameter PMA_REG_ALG_CTLE_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_CTLE_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_CTLE_INITDAC_6 = 0,
    parameter PMA_REG_ALG_CTLE_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_2_0 = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_4_3 = 2,
    parameter PMA_REG_ALG_CTLEOFS_FLIPDIR_I = "TRUE",
    parameter PMA_REG_ALG_CTLEOFS_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_3_0 = 0,
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_6_4 = 4,
    parameter PMA_REG_ALG_CTLEOFS_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_SHIFT_I = 4,
    parameter PMA_REG_ALG_DFE_CTLE_PWD = "FALSE",
    parameter PMA_REG_ALG_H1_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H1_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_H1_INITDAC_6 = 0,
    parameter PMA_REG_ALG_H1_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_SHIFT_I = 4,
    parameter PMA_REG_ALG_H2_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H2_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H2_INITDAC_5_1 = 0,
    parameter PMA_REG_ALG_H2_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_SHIFT_I_1_0 = 0,
    parameter integer PMA_REG_ALG_H2_SHIFT_I_2 = 1,
    parameter PMA_REG_ALG_H3_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H3_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_INITDAC_4_0 = 0,
    parameter integer PMA_REG_ALG_H3_INITDAC_5 = 1,
    parameter PMA_REG_ALG_H3_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_SHIFT_I = 4,
    parameter PMA_REG_ALG_H4_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H4_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H4_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_H4_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_SHIFT_I = 4,
    parameter PMA_REG_ALG_H5_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H5_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_INITDAC = 16,
    parameter PMA_REG_ALG_H5_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_SHIFT_I = 4,
    parameter PMA_REG_ALG_H6_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H6_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_H6_INITDAC_4_3 = 2,
    parameter PMA_REG_ALG_H6_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_HCTLE_OFS_1_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OFS_3_2 = 2,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_6 = 1,
    parameter PMA_REG_ALG_HCTLE_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQH_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQH_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_REG_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_LEQL_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQL_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQL_REG_PRESELECT_I = 7,
    parameter integer PMA_REG_ALG_LEQL_REG_SHIFT_I = 4,
    parameter PMA_REG_ALG_NEXTBIT_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_6_0 = 127,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_14_7 = 255,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_19_15 = 31,
    parameter integer PMA_REG_ALG_SOFS_DACWIN_I = 1,
    parameter PMA_REG_ALG_SOFS_FLIP_DIR_I = "TRUE",
    parameter PMA_REG_ALG_SOFS_FORCE_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_5_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_6 = 1,
    parameter integer PMA_REG_ALG_SOFS_FORCENUM_I = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_6_3 = 8,
    parameter integer PMA_REG_ALG_SOFS_SHIFT_I = 1,
    parameter PMA_REG_ALG_SOFS_SKIP_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0 = 254,
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8 = 15,
    parameter PMA_REG_ALG_ST_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_ST_FORCEN = "FALSE",
    parameter PMA_REG_ALG_ST_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_ST_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_ST_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_ST_RECALEN = "FALSE",
    parameter integer PMA_REG_ALG_ST_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_ST_STARTCNT_7_0 = 0,
    parameter integer PMA_REG_ALG_ST_STARTCNT_15_8 = 128,
    parameter integer PMA_REG_ALG_ST_STARTCNT_19_16 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_3_0 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_11_4 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_17_12 = 2,
    parameter integer PMA_REG_ALG_ST_TOPTAP_1_0 = 3,
    parameter integer PMA_REG_ALG_ST_TOPTAP_3_2 = 3,
    parameter integer PMA_REG_ALG_SWCLK_DIV = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_3_0 = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_4 = 1,
    parameter integer PMA_REG_ALG_TAPA_NUM = 7,
    parameter integer PMA_REG_ALG_TAPB_DAC_0 = 0,
    parameter integer PMA_REG_ALG_TAPB_DAC_4_1 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_3_0 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_5_4 = 0,
    parameter integer PMA_REG_ALG_TAPC_DAC = 16,
    parameter integer PMA_REG_ALG_TAPC_NUM_0 = 1,
    parameter integer PMA_REG_ALG_TAPC_NUM_5_1 = 4,
    parameter integer PMA_REG_ALG_TAPD_DAC_2_0 = 0,
    parameter integer PMA_REG_ALG_TAPD_DAC_4_3 = 2,
    parameter integer PMA_REG_ALG_TAPD_NUM = 10,
    parameter PMA_REG_ALG_VP_FLIPDIR_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_GRN_SHIFT_I = 5,
    parameter PMA_REG_ALG_VP_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_IDEAL_2_0 = 0,
    parameter integer PMA_REG_ALG_VP_IDEAL_6_3 = 10,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_3_0 = 0,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_6_4 = 0,
    parameter PMA_REG_ALG_VP_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_VP_RED_SHIFT_I = 5,
    parameter integer PMA_REG_ALG_VPOFS_SEL_0 = 0,
    parameter integer PMA_REG_ALG_VPOFS_SEL_2_1 = 1,
    parameter integer PMA_REG_ALG_H1_UPBOUND_5_0 = 55,
    parameter integer PMA_REG_ALG_H1_UPBOUND_6 = 1,
    parameter PMA_REG_ALG_CTLEOFS_PWDN = "FALSE",
    parameter PMA_REG_ALG_LEQH_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_AGC_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_AGC_INITDAC = 10,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_1_0 = 3,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_3_2 = 0,
    parameter PMA_REG_ALG_AGC_OVERWREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_PWD = "FALSE",
    parameter integer PMA_REG_ALG_AGC_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_0 = 1,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_3_1 = 7,
    parameter integer PMA_REG_ALG_AGC_WAITSEL = 11,
    parameter PMA_REG_PI_CTRL_SEL_RX = "FALSE",
    parameter integer PMA_REG_PI_CTRL_RX_4_0 = 0,
    parameter integer PMA_REG_PI_CTRL_RX_7_5 = 0,
    parameter PMA_CFG_RX_LANE_POWERUP = "ON",
    parameter PMA_CFG_RX_PMA_RSTN = "TRUE",
    parameter PMA_INT_PMA_RX_MASK_0 = "FALSE",
    parameter PMA_INT_PMA_RX_CLR_0 = "FALSE",
    parameter PMA_CFG_CTLE_ADP_RSTN = "TRUE",
    parameter PMA_CFG_RX_CDR_RSTN = "TRUE",
    parameter PMA_CFG_RX_CLKPATH_RSTN = "TRUE",
    parameter PMA_CFG_RX_DFE_RSTN = "TRUE",
    parameter PMA_CFG_RX_LEQ_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIDING_RSTN = "TRUE",
    parameter PMA_CFG_RX_EYE_RSTN = "TRUE",
    parameter PMA_CFG_RX_CTLE_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLICER_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIP_RSTN = "TRUE",
    parameter integer PMA_REG_TX_BEACON_TIMER_SEL = 0,
    parameter PMA_REG_TX_BIT_CONV = "FALSE",
    parameter integer PMA_REG_TX_RES_CAL = 50,
    parameter integer PMA_REG_TX_UDP_DATA_20 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_26_21 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_34_27 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_39_25 = 0,
    parameter integer PMA_REG_TX_BUSWIDTH_EN = 0,
    parameter PMA_REG_TX_PD_POST = "OFF",
    parameter PMA_REG_TX_PD_POST_OW = "FALSE",
    parameter PMA_REG_TX_BUSWIDTH = "20BIT",
    parameter integer PMA_REG_EI_PCLK_DELAY_SEL = 0,
    parameter integer PMA_REG_TX_AMP_DAC0 = 25,
    parameter integer PMA_REG_TX_AMP_DAC1 = 19,
    parameter integer PMA_REG_TX_AMP_DAC2 = 14,
    parameter integer PMA_REG_TX_AMP_DAC3 = 9,
    parameter PMA_REG_TX_RXDET_THRESHOLD = "84MV",
    parameter PMA_REG_TX_BEACON_OSC_CTRL = "FALSE",
    parameter integer PMA_REG_TX_PRBS_GEN_WIDTH_SEL = 0,
    parameter PMA_REG_TX_TX2RX_SLPBACK_EN = "FALSE",
    parameter PMA_REG_TX_PCLK_EDGE_SEL = "FALSE",
    parameter PMA_REG_TX_PRBS_GEN_EN = "FALSE",
    parameter PMA_REG_TX_PRBS_SEL = "PRBS7",
    parameter integer PMA_REG_TX_UDP_DATA_7_TO_0 = 5,
    parameter integer PMA_REG_TX_UDP_DATA_15_TO_8 = 235,
    parameter integer PMA_REG_TX_UDP_DATA_19_TO_16 = 3,
    parameter integer PMA_REG_TX_FIFO_WP_CTRL = 4,
    parameter PMA_REG_TX_FIFO_EN = "FALSE",
    parameter integer PMA_REG_TX_DATA_MUX_SEL = 0,
    parameter PMA_REG_TX_ERR_INSERT = "FALSE",
    parameter PMA_REG_TX_SATA_EN = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON_OW = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON = "TRUE",
    parameter integer PMA_REG_TX_CFG_POST1 = 0,
    parameter integer PMA_REG_TX_CFG_POST2 = 0,
    parameter integer PMA_REG_TX_OOB_DELAY_SEL = 0,
    parameter PMA_REG_TX_POLARITY = "NORMAL",
    parameter PMA_REG_TX_LS_MODE_EN = "FALSE",
    parameter PMA_REG_RX_JTAG_OE = "TRUE",
    parameter integer PMA_REG_RX_ACJTAG_VHYSTSEL = 0,
    parameter PMA_REG_TX_RES_CAL_EN = "FALSE",
    parameter integer PMA_REG_RX_TERM_MODE_CTRL = 5,
    parameter PMA_REG_PLPBK_TXPCLK_EN = "FALSE",
    parameter integer PMA_REG_CLK_SEL_STROBE_TXPCLK = 2,
    parameter integer PMA_REG_TX_PH_SEL_0 = 1,
    parameter integer PMA_REG_TX_PH_SEL_6_1 = 0,
    parameter integer PMA_REG_TX_CFG_PRE = 0,
    parameter integer PMA_REG_TX_CFG_MAIN = 0,
    parameter integer PMA_REG_CFG_POST = 0,
    parameter PMA_REG_PD_MAIN = "TRUE",
    parameter PMA_REG_PD_PRE = "TRUE",
    parameter integer PMA_REG_TX_RXDET_TIMER_SEL = 87,
    parameter PMA_REG_TX_PI_CUR_BUF = "10GHz",
    parameter PMA_REG_TX_MOD_STAND_BY_EN = "FALSE",
    parameter PMA_REG_STATE_STAND_BY_SEL = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_POLAR_CTRL = "FALSE",
    parameter PMA_REG_TX_FREERUN_PD = "TRUE",
    parameter PMA_REG_TX_CHANGE_ON_SEL = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_CTRL = "FALSE",
    parameter integer PMA_REG_TX_FREERUN_RATE_0 = 0,
    parameter integer PMA_REG_TX_FREERUN_RATE_1 = 0,
    parameter PMA_REG_TX_FREERUN_RATE_OW = "FALSE",
    parameter PMA_REG_TX_RST_SYNC_CLK_SEL = "TRUE",
    parameter integer PMA_REG_TX_PI_CTRL_SEL = 0,
    parameter integer PMA_REG_TX_PI_CTRL = 0,
    parameter PMA_LANE_POWERUP = "TRUE",
    parameter PMA_POR_N = "TRUE",
    parameter PMA_TX_LANE_POWERUP = "TRUE",
    parameter PMA_TX_PMA_RSTN = "TRUE",
    parameter PMA_LPLL_POWERUP = "TRUE",
    parameter PMA_LPLL_RSTN = "TRUE",
    parameter PMA_LPLL_LOCKDET_RSTN = "TRUE",
    parameter integer PMA_REG_LPLL_PFDDELAY_SEL = 1,
    parameter PMA_REG_LPLL_PFDDELAY_EN = "TRUE",
    parameter integer PMA_REG_LPLL_VCTRL_SET = 0,
    parameter PMA_LPLL_CHARGE_PUMP_CTRL = "type",
    parameter PMA_LPLL_REFDIV = "DIV1",
    parameter integer PMA_LPLL_FBDIV = 38,
    parameter integer PMA_LPLL_LPF_RES = 1,
    parameter integer PMA_LPLL_REFLOSS_READY = 0,
    parameter integer PMA_LPLL_LOCKED_PFDDELAY = 0,
    parameter integer PMA_LPLL_MCLK_SEL = 0,
    parameter integer PMA_LPLL_TEST_SEL = 0,
    parameter PMA_LPLL_TEST_SIG_HALF_EN = "TRUE",
    parameter PMA_LPLL_TEST_V_EN = "FALSE",
    parameter PMA_LPLL_MCLK_EN = "TRUE",
    parameter integer PMA_LPLL_MCLK_DET_CTL = 16,
    parameter integer PMA_LPLL_LOCKDET_REFCT = 3,
    parameter integer PMA_LPLL_LOCKDET_FBCT = 3,
    parameter integer PMA_LPLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_LPLL_LOCKDET_ITER = 1,
    parameter integer PMA_LPLL_UNLOCKDET_ITER = 2,
    parameter integer PMA_LPLL_LOCKDET_EN_OW = 0,
    parameter integer PMA_LPLL_LOCKDET_EN = 0,
    parameter integer PMA_LPLL_LOCKDET_MODE = 0,
    parameter integer PMA_LPLL_LOCKDET_OW = 0,
    parameter integer PMA_LPLL_LOCKDETED = 0,
    parameter integer PMA_LPLL_UNLOCKDET_OW = 0,
    parameter integer PMA_LPLL_UNLOCKDETED = 0,
    parameter integer PMA_LPLL_LOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_UNLOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_LOCKDET_REPEAT = 0,
    parameter integer PMA_LPLL_NOFBCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_NOREFCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_READY_OR_LOCK = 0,
    parameter integer PMA_LPLL_READY = 0,
    parameter integer PMA_LPLL_READY_OW = 0,
    parameter PMA_REG_TXCLK_SEL = "HPLL",
    parameter PMA_REG_RXCLK_SEL = "HPLL",
    parameter integer PMA_REG_TEST_BUF = 0,
    parameter PMA_REG_RX_DEF_SEL0 = "18.75uA",
    parameter PMA_REG_RX_DEF_SEL1 = "18.75uA",
    parameter PMA_REG_TX_DIV_SEL = "25uA",
    parameter PMA_REG_LPLL_AMP_SEL = "25uA",
    parameter PMA_REG_LPLL_VCO_SEL = "25uA",
    parameter PMA_REG_LPLL_CHARGE_PUMP_SEL = "25uA",
    parameter PMA_REG_RX_EQ0_SEL = "56.25uA",
    parameter PMA_REG_RX_EQ1_SEL = "56.25uA",
    parameter PMA_REG_RX_PGA_SEL = "56.25uA",
    parameter integer PMA_REG_CHL_TEST = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_7_0 = 255,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_15_8 = 247,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_18_16 = 7,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_21_19 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_29_22 = 0,
    parameter integer PMA_REG_IBIAS_STATIC_SEL_37_30 = 1,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_7_0 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_15_8 = 0,
    parameter integer PMA_REG_IBIAS_DYNAMIC_PD_18_16 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_4_0 = 31,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_8_5 = 15,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_12_9 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_SEL_17_13 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_2_0 = 0,
    parameter integer PMA_REG_IBIAS_STA_CUR_PD_8_3 = 0,
    parameter PMA_REG_BANDGAP_VOL_SEL = "BANDGAP",
    parameter integer PMA_REG_BANDGAP_TEST = 0
) (
    output P_CFG_READY,
    output [7:0] P_CFG_RDATA,
    output P_CFG_INT,
    output [24:0] LANE_COUT_BUS_FORWARD,
    output [1:0] LANE_COUT_BUS_BACKWARD,
    output P_RX_PRBS_ERROR,
    output P_PCS_RX_MCB_STATUS,
    output P_PCS_LSM_SYNCED,
    output [87:0] P_RDATA,
    output P_RXDVLD,
    output P_RXDVLD_H,
    output [5:0] P_RXSTATUS,
    output [2:0] P_EM_ERROR_CNT,
    output P_LPLL_READY,
    output P_RX_SIGDET_STATUS,
    output P_RX_SATA_COMINIT,
    output P_RX_SATA_COMWAKE,
    output P_RX_LS_DATA,
    output P_RX_READY,
    output [19:0] P_TEST_STATUS,
    output P_TX_RXDET_STATUS,
    output P_RCLK2FABRIC,
    output P_TCLK2FABRIC,
    output P_CA_ALIGN_RX,
    output P_CA_ALIGN_TX,
    output P_TX_SDN,
    output P_TX_SDP,
    input P_RX_CLK_FR_CORE,
    input P_RCLK2_FR_CORE,
    input P_TX_CLK_FR_CORE,
    input P_TCLK2_FR_CORE,
    input P_PCS_RX_RST,
    input P_PCS_TX_RST,
    input P_EXT_BRIDGE_PCS_RST,
    input P_CFG_RST,
    input P_CFG_CLK,
    input P_CFG_PSEL,
    input P_CFG_ENABLE,
    input P_CFG_WRITE,
    input [11:0] P_CFG_ADDR,
    input [7:0] P_CFG_WDATA,
    input [24:0] LANE_CIN_BUS_FORWARD,
    input [1:0] LANE_CIN_BUS_BACKWARD,
    input [87:0] P_TDATA,
    input P_PCIE_EI_H,
    input P_PCIE_EI_L,
    input [15:0] P_TX_DEEMP,
    input [1:0] P_TX_DEEMP_POST_SEL,
    input P_BLK_ALIGN_CTRL,
    input P_TX_ENC_TYPE,
    input P_RX_DEC_TYPE,
    input P_PCS_BIT_SLIP,
    input P_PCS_WORD_ALIGN_EN,
    input P_RX_POLARITY_INVERT,
    input P_PCS_MCB_EXT_EN,
    input P_PCS_NEAREND_LOOP,
    input P_PCS_FAREND_LOOP,
    input P_PMA_NEAREND_PLOOP,
    input P_PMA_NEAREND_SLOOP,
    input P_PMA_FAREND_PLOOP,
    input P_PCS_PRBS_EN,
    input P_LANE_POWERDOWN,
    input P_LANE_RST,
    input P_RX_LANE_POWERDOWN,
    input P_RX_PMA_RST,
    input P_RX_CDR_RST,
    input P_RX_CLKPATH_RST,
    input P_RX_DFE_RST,
    input P_RX_LEQ_RST,
    input P_RX_SLIDING_RST,
    input P_RX_DFE_EN,
    input P_RX_T1_EN,
    input P_RX_CDRX_EN,
    input P_RX_T1_DFE_EN,
    input P_RX_T2_DFE_EN,
    input P_RX_T3_DFE_EN,
    input P_RX_T4_DFE_EN,
    input P_RX_T5_DFE_EN,
    input P_RX_T6_DFE_EN,
    input P_RX_SLIDING_EN,
    input P_RX_EYE_RST,
    input P_RX_EYE_EN,
    input [7:0] P_RX_EYE_TAP,
    input [7:0] P_RX_PIC_EYE,
    input [7:0] P_RX_PIC_FASTLOCK,
    input P_RX_PIC_FASTLOCK_STROBE,
    input P_EM_RD_TRIGGER,
    input [1:0] P_EM_MODE_CTRL,
    input P_RX_CTLE_DCCAL_RST,
    input P_RX_SLICER_DCCAL_RST,
    input P_RX_SLICER_DCCAL_EN,
    input P_RX_CTLE_DCCAL_EN,
    input P_RX_SLIP_RST,
    input P_RX_SLIP_EN,
    input P_LPLL_POWERDOWN,
    input P_LPLL_RST,
    input P_LPLL_LOCKDET_RST,
    input P_TX_LS_DATA,
    input P_TX_BEACON_EN,
    input P_TX_SWING,
    input P_TX_RXDET_REQ,
    input [1:0] P_TX_RATE,
    input [2:0] P_TX_BUSWIDTH,
    input [2:0] P_TX_FREERUN_BUSWIDTH,
    input [2:0] P_TX_MARGIN,
    input P_TX_PMA_RST,
    input P_TX_LANE_POWERDOWN,
    input P_TX_PIC_EN,
    input [1:0] P_RX_RATE,
    input [2:0] P_RX_BUSWIDTH,
    input P_RX_HIGHZ,
    input [7:0] P_CIM_CLK_ALIGNER_RX,
    input [7:0] P_CIM_CLK_ALIGNER_TX,
    input P_ALIGN_MODE_VALID_RX,
    input [1:0] P_ALIGN_MODE_RX,
    input P_ALIGN_MODE_VALID_TX,
    input [2:0] P_ALIGN_MODE_TX,
    input PMA_HPLL_CK0,
    input PMA_HPLL_CK90,
    input PMA_HPLL_CK180,
    input PMA_HPLL_CK270,
    input PMA_HPLL_READY_IN,
    input PMA_HPLL_REFCLK_IN,
    input PMA_TX_SYNC_HPLL_IN,
    input P_LPLL_REFCLK_IN,
    input P_TX_RATE_CHANGE_ON_0,
    input P_TX_RATE_CHANGE_ON_1,
    input P_TX_SYNC,
    input P_RX_SDN,
    input P_RX_SDP,
    input P_CDR_PICTRL_OW,
    input [7:0] P_CDR_PICTRL_OW_VAL
)  ;
endmodule


module GTP_HSSTHP_LANE_t
#(
    parameter PCS_DYN_DLY_SEL_RX = "FALSE",
    parameter PCS_PMA_RCLK_POLINV = "PMA_RCLK",
    parameter PCS_PCS_RCLK_SEL = "RCLK",
    parameter PCS_GEAR_RCLK_SEL = "RCLK",
    parameter PCS_RCLK2FABRIC_SEL = "HARD_1",
    parameter PCS_SCAN_INTERVAL_RX = "4_CLOCKS",
    parameter PCS_BRIDGE_RCLK_SEL = "RCLK",
    parameter PCS_RCLK_POLINV = "RCLK",
    parameter PCS_TO_FABRIC_CLK_SEL = "PMA_RCLK",
    parameter PCS_CLK2ALIGNER_SEL = "TO_FABRIC_CLK",
    parameter PCS_TO_FABRIC_CLK_DIV_EN = "FALSE",
    parameter PCS_AUTO_NEAR_LOOP_EN = "FALSE",
    parameter PCS_PCS_RCLK_EN = "FALSE",
    parameter PCS_BRIDGE_PCS_RCLK_EN_SEL = "HARD_1",
    parameter PCS_BRIDGE_RCLK_EN_SEL = "HARD_0",
    parameter PCS_GEAR_RCLK_EN_SEL = "HARD_0",
    parameter PCS_NEGEDGE_EN_RX = "FALSE",
    parameter PCS_PCS_RX_RSTN = "FALSE",
    parameter PCS_BRIDGE_PCS_RSTN = "FALSE",
    parameter PCS_TO_FABRIC_RST_EN = "FALSE",
    parameter PCS_BYPASS_GEAR_RRSTN = "FALSE",
    parameter PCS_BYPASS_BRIDGE_RRSTN = "FALSE",
    parameter PCS_ALIGNER_EN_RX = "FALSE",
    parameter PCS_RX_SLAVE = "MASTER",
    parameter integer PCS_RX_CA = 0,
    parameter integer PCS_SUM_THRESHOLD_RX = 0,
    parameter integer PCS_AVG_CYCLES_RX = 0,
    parameter PCS_REG_PMA_RX2TX_PLOOP_EN = "FALSE",
    parameter PCS_REG_PMA_RX2TX_PLOOP_FIFOEN = "FALSE",
    parameter integer PCS_STEP_SIZE_RX = 0,
    parameter integer PCS_REV_CNT_LIMIT_RX = 0,
    parameter integer PCS_FILTER_CNT_SIZE_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_3_0 = 0,
    parameter integer PCS_DLY_REC_SIZE_RX = 0,
    parameter integer PCS_ALIGN_THRD_RX = 0,
    parameter integer PCS_DLY_ADJUST_SIZE_RX_4 = 0,
    parameter PCS_CFG_DEC_TYPE_EN = "FALSE",
    parameter PCS_RXBRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_GE_AUTO_EN = "FALSE",
    parameter PCS_RXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_RXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_IFG_EN = "FALSE",
    parameter PCS_FLP_FULL_CHK_EN = "FALSE",
    parameter PCS_FLP_EMPTY_CHK_EN = "FALSE",
    parameter PCS_RX_POLARITY_INV = "DELAY",
    parameter PCS_FARLP_PWR_REDUCTION = "FALSE",
    parameter PCS_RXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_WDALIGN_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXDEC_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_RXTEST_PWR_REDUCTION = "NORMAL",
    parameter integer PCS_WA_SOS_DET_TOL = 0,
    parameter integer PCS_WA_SE_DET_TOL = 0,
    parameter PCS_RX_SAMPLE_UNION = "FALSE",
    parameter PCS_NEAR_LOOP = "FALSE",
    parameter PCS_BYPASS_WORD_ALIGN = "FALSE",
    parameter PCS_BYPASS_DENC = "FALSE",
    parameter PCS_RX_ERRCNT_CLR = "FALSE",
    parameter PCS_RX_CODE_MODE = "DUAL_8B10B",
    parameter PCS_RX_BYPASS_GEAR = "FALSE",
    parameter PCS_ERRDETECT_SILENCE = "FALSE",
    parameter PCS_RX_DATA_MODE = "8BIT",
    parameter PCS_CA_DYN_CLY_EN_RX = "FALSE",
    parameter PCS_CFG_APATTERN_STATUS_DELAY = "DELAY_ONE_CYCLE",
    parameter PCS_RX_PRBS_MODE = "DISABLE",
    parameter PCS_ALIGN_MODE = "1GB",
    parameter PCS_COMMA_DET_MODE = "PATTERN_DETECT",
    parameter integer PCS_RAPID_VMIN_1 = 0,
    parameter integer PCS_RAPID_VMIN_2 = 0,
    parameter PCS_RXBU_WIDER_EN = "40/20BIT",
    parameter integer PCS_RAPID_IMAX = 0,
    parameter PCS_RX_SPLIT = "SPLIT_22BIT_11BIT",
    parameter integer PCS_RXBRG_END_PACKET_9_8 = 0,
    parameter integer PCS_RXBRG_END_PACKET_7_0 = 0,
    parameter integer PCS_CTC_MAX_DEL = 0,
    parameter integer PCS_COMMA_REG0_9_8 = 0,
    parameter integer PCS_COMMA_REG1_9_8 = 0,
    parameter integer PCS_COMMA_MASK_9_8 = 0,
    parameter integer PCS_COMMA_REG0_7_0 = 0,
    parameter integer PCS_COMMA_REG1_7_0 = 0,
    parameter integer PCS_COMMA_MASK_7_0 = 0,
    parameter integer PCS_FLP_WRADDR_START = 0,
    parameter integer PCS_FLP_RDADDR_START = 0,
    parameter PCS_CFG_RX_BRIDGE_CLK_POLINV = "FALSE",
    parameter PCS_CTC_MODE_RD_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AFULL = 0,
    parameter PCS_FAST_LOCK_GEAR_EN = "FALSE",
    parameter PCS_CTC_MODE_WR_SEL = "NOMINAL_EMPTY",
    parameter integer PCS_CTC_AEMPTY = 0,
    parameter PCS_CTC_MODE = "ONE_BYTE",
    parameter PCS_RXBRIDGE_MODE = "BYPASS",
    parameter integer PCS_CTC_ADD_MAX = 0,
    parameter PCS_CFG_PHDET_EN_RX = "FALSE",
    parameter integer PCS_WA_SDS_DET_TOL = 0,
    parameter PCS_CEB_MODE = "10GB",
    parameter PCS_APATTERN_MODE = "ONE_BYTE",
    parameter PCS_A_REG0_8 = "FALSE",
    parameter integer PCS_RXBRG_WADDR_START = 0,
    parameter PCS_A_REG1_8 = "FALSE",
    parameter integer PCS_RXBRG_RADDR_START = 0,
    parameter integer PCS_A_REG0_7_0 = 0,
    parameter integer PCS_A_REG1_7_0 = 0,
    parameter integer PCS_CEB_RAPIDLS_MMAX = 0,
    parameter integer PCS_CEB_DETECT_TIME = 0,
    parameter integer PCS_WL_FIFO_RD = 0,
    parameter integer PCS_SKIP_REG0_9_8 = 0,
    parameter integer PCS_SKIP_REG0_7_0 = 0,
    parameter integer PCS_CFG_CONTI_SKP_SET = 0,
    parameter PCS_CFG_RX_BASE_ADV_MODE = "BASE_MODE",
    parameter integer PCS_SKIP_REG1_9_8 = 0,
    parameter integer PCS_SKIP_REG2_9_8 = 0,
    parameter integer PCS_SKIP_REG3_9_8 = 0,
    parameter integer PCS_SKIP_REG1_7_0 = 0,
    parameter integer PCS_SKIP_REG2_7_0 = 0,
    parameter integer PCS_SKIP_REG3_7_0 = 0,
    parameter integer PCS_CFG_PRBS_ERR_O_SEL = 0,
    parameter integer PCS_CFG_PD_DELAY_RX = 0,
    parameter integer PCS_WR_START_GAP = 0,
    parameter integer PCS_MIN_IFG = 0,
    parameter PCS_INT_RX_MASK_0 = "FALSE",
    parameter PCS_INT_RX_MASK_1 = "FALSE",
    parameter PCS_INT_RX_MASK_2 = "FALSE",
    parameter PCS_INT_RX_MASK_3 = "FALSE",
    parameter PCS_INT_RX_MASK_4 = "FALSE",
    parameter PCS_INT_RX_MASK_5 = "FALSE",
    parameter PCS_INT_RX_CLR_5 = "FALSE",
    parameter PCS_INT_RX_CLR_4 = "FALSE",
    parameter PCS_INT_RX_CLR_3 = "FALSE",
    parameter PCS_INT_RX_CLR_2 = "FALSE",
    parameter PCS_INT_RX_CLR_1 = "FALSE",
    parameter PCS_INT_RX_CLR_0 = "FALSE",
    parameter PCS_EM_CNT_RD_EN = "FALSE",
    parameter PCS_EM_CTRL_SEL = "SIGNAL_CTRL",
    parameter PCS_EM_MODE_CTRL = "HOLD",
    parameter PCS_EM_RD_CONDITION = "TRIGGER",
    parameter integer PCS_EM_SP_PATTERN_7_0 = 0,
    parameter integer PCS_EM_SP_PATTERN_15_8 = 0,
    parameter integer PCS_EM_SP_PATTERN_23_16 = 0,
    parameter integer PCS_EM_SP_PATTERN_31_24 = 0,
    parameter integer PCS_EM_SP_PATTERN_39_32 = 0,
    parameter integer PCS_EM_SP_PATTERN_47_40 = 0,
    parameter integer PCS_EM_SP_PATTERN_55_48 = 0,
    parameter integer PCS_EM_SP_PATTERN_63_56 = 0,
    parameter integer PCS_EM_SP_PATTERN_71_64 = 0,
    parameter integer PCS_EM_SP_PATTERN_79_72 = 0,
    parameter integer PCS_EM_PMA_MASK_7_0 = 0,
    parameter integer PCS_EM_PMA_MASK_15_8 = 0,
    parameter integer PCS_EM_PMA_MASK_23_16 = 0,
    parameter integer PCS_EM_PMA_MASK_31_24 = 0,
    parameter integer PCS_EM_PMA_MASK_39_32 = 0,
    parameter integer PCS_EM_PMA_MASK_47_40 = 0,
    parameter integer PCS_EM_PMA_MASK_55_48 = 0,
    parameter integer PCS_EM_PMA_MASK_63_56 = 0,
    parameter integer PCS_EM_PMA_MASK_71_64 = 0,
    parameter integer PCS_EM_PMA_MASK_79_72 = 0,
    parameter integer PCS_EM_EYED_MASK_7_0 = 0,
    parameter integer PCS_EM_EYED_MASK_15_8 = 0,
    parameter integer PCS_EM_EYED_MASK_23_16 = 0,
    parameter integer PCS_EM_EYED_MASK_31_24 = 0,
    parameter integer PCS_EM_EYED_MASK_39_32 = 0,
    parameter integer PCS_EM_EYED_MASK_47_40 = 0,
    parameter integer PCS_EM_EYED_MASK_55_48 = 0,
    parameter integer PCS_EM_EYED_MASK_63_56 = 0,
    parameter integer PCS_EM_EYED_MASK_71_64 = 0,
    parameter integer PCS_EM_EYED_MASK_79_72 = 0,
    parameter integer PCS_EM_PRESCALE = 0,
    parameter PCS_CFG_TEST_STATUS_SEL = "SEL_PMA_TEST_STATUS_INT",
    parameter integer PCS_CFG_DIFF_CNT_BND_RX = 0,
    parameter PCS_CFG_FLT_SEL_RX = "FALSE",
    parameter integer PCS_FILTER_BND_RX = 0,
    parameter PCS_TCLK2FABRIC_DIV_RST_M = "FALSE",
    parameter PCS_TX_PMA_TCLK_POLINV = "PMA_TCLK",
    parameter PCS_TX_TCLK_POLINV = "TCLK",
    parameter PCS_PCS_TCLK_SEL = "PMA_TCLK",
    parameter PCS_GEAR_TCLK_SEL = "PMA_TCLK",
    parameter PCS_TX_BRIDGE_TCLK_SEL = "TCLK",
    parameter PCS_TCLK2ALIGNER_SEL = "PMA_TCLK",
    parameter CA_DYN_DLY_EN_TX = "FALSE",
    parameter PCS_TX_PCS_CLK_EN_SEL = "HARDWIRED1",
    parameter PCS_TX_GEAR_CLK_EN_SEL = "HARDWIRED0",
    parameter PCS_TCLK2FABRIC_DIV_EN = "FALSE",
    parameter PCS_TCLK2FABRIC_SEL = "CLK2ALIGNER_N_DIV2",
    parameter integer DLY_ADJUST_SIZE_TX = 0,
    parameter PCS_TX_PCS_TX_RSTN = "FALSE",
    parameter PCS_TX_CA_RSTN = "FALSE",
    parameter PCS_TX_SLAVE = "MASTER",
    parameter integer PCS_TX_CA = 0,
    parameter integer PCS_CFG_PI_CLK_SEL = 0,
    parameter PCS_CFG_PI_CLK_EN_SEL = "CLK_EN_ALWAYS1",
    parameter integer PCS_CFG_PI_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_SUM_THRESHOLD_TX = 0,
    parameter integer PCS_CFG_AVG_CYCLES_TX = 0,
    parameter PCS_CFG_NEGEDGE_EN_TX = "FALSE",
    parameter integer PCS_CFG_ALIGN_THRD_TX = 0,
    parameter integer PCS_CFG_SCAN_INTERVAL_TX = 0,
    parameter integer PCS_CFG_STEP_SIZE_TX = 0,
    parameter integer PCS_CFG_REV_CNT_LIMIT_TX = 0,
    parameter integer PCS_CFG_FILTER_CNT_SIZE_TX = 0,
    parameter integer PCS_CFG_PI_DEFAULT_TX = 0,
    parameter PCS_CFG_PHDET_EN_TX = "FALSE",
    parameter PCS_PMA_TX2RX_PLOOP_EN = "FALSE",
    parameter PCS_PMA_TX2RX_SLOOP_EN = "FALSE",
    parameter PCS_CFG_DYN_DLY_SEL_TX = "FALSE",
    parameter integer PCS_CFG_DLY_REC_SIZE_TX = 0,
    parameter PCS_TX_DATA_WIDTH_MODE = "8BIT",
    parameter PCS_TX_BYPASS_BRIDGE_UINT = "FALSE",
    parameter PCS_TX_BYPASS_BRIDGE_FIFO = "FALSE",
    parameter PCS_TX_BYPASS_GEAR = "FALSE",
    parameter PCS_TX_BYPASS_ENC = "FALSE",
    parameter PCS_TX_BYPASS_BIT_SLIP = "FALSE",
    parameter PCS_TX_BRIDGE_GEAR_SEL = "FALSE",
    parameter PCS_TXBRG_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXGEAR_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXENC_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBSLP_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXPRBS_PWR_REDUCTION = "NORMAL",
    parameter PCS_TXBRG_FULL_CHK_EN = "FALSE",
    parameter PCS_TXBRG_EMPTY_CHK_EN = "FALSE",
    parameter PCS_TX_ENCODER_MODE = "DUAL_8B10B",
    parameter PCS_TX_PRBS_MODE = "DISABLE",
    parameter PCS_TX_DRIVE_REG_MODE = "NO_CHANGE",
    parameter integer PCS_TX_BIT_SLIP_CYCLES = 0,
    parameter PCS_TX_BASE_ADV_MODE = "BASE",
    parameter PCS_TX_GEAR_SPLIT = "NO_SPILT",
    parameter PCS_RX_BRIDGE_CLK_POLINV = "N_CLK_INVERT",
    parameter PCS_PRBS_ERR_LPBK = "FALSE",
    parameter PCS_TX_INSERT_ER = "FALSE",
    parameter PCS_ENABLE_PRBS_GEN = "FALSE",
    parameter PCS_FAR_LOOP = "FALSE",
    parameter PCS_CFG_ENC_TYPE_EN = "FALSE",
    parameter integer PCS_TXBRG_WADDR_START = 0,
    parameter integer PCS_TXBRG_RADDR_START = 0,
    parameter PCS_CFG_TX_PIC_EN = "DISABLE",
    parameter PCS_CFG_PIC_DIRECT_INV = "FALSE",
    parameter PCS_CFG_PI_MOD_CLK_EN = "FALSE",
    parameter PCS_CFG_TX_MODULATOR_OW_EN = "FALSE",
    parameter PCS_CFG_TX_PI_SSC_MODE_EN = "FALSE",
    parameter PCS_CFG_TX_PI_OFFSET_MODE_EN = "FALSE",
    parameter integer PCS_CFG_TX_PI_SSC_MODE_SEL = 0,
    parameter PCS_CFG_TXDEEMPH_EN = "FALSE",
    parameter PCS_PI_STROBE_SEL = "FALSE",
    parameter PCS_CFG_TX_PIC_GREY_SEL = "FALSE",
    parameter PCS_CFG_PIC_RENEW_INV = "NORMAL",
    parameter integer PCS_CFG_NUM_PIC = 0,
    parameter PCS_CFG_TXPIC_OW_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_OW_VALUE_0_7 = 0,
    parameter PCS_INT_TX_MASK_0 = "FALSE",
    parameter PCS_INT_TX_MASK_1 = "FALSE",
    parameter PCS_INT_TX_MASK_2 = "FALSE",
    parameter PCS_TX_WPTR_SEL = "FALSE",
    parameter PCS_INT_TX_CLR_2 = "FALSE",
    parameter PCS_INT_TX_CLR_1 = "FALSE",
    parameter PCS_INT_TX_CLR_0 = "FALSE",
    parameter integer PCS_CFG_PD_DELAY_TX = 0,
    parameter integer PCS_CFG_DIFF_CNT_BND_TX = 0,
    parameter PCS_CFG_PD_CLK_FR_CORE_SEL = "FALSE",
    parameter PCS_CFG_FLT_SEL_TX = "FALSE",
    parameter integer PCS_FILTER_BND_TX = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_7_0 = 0,
    parameter PCS_CFG_TX_SSC_MODULATOR_EN = "FALSE",
    parameter integer PCS_CFG_TX_SSC_SCALE2_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_SCALE_SEL = 0,
    parameter integer PCS_CFG_TX_SSC_RANGE_8_9 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_7_0 = 0,
    parameter integer PCS_CFG_TX_SSC_MODULATION_STEP_8 = 0,
    parameter integer PCS_CFG_TX_SSC_OFFSET_8_9 = 0,
    parameter PMA_REG_CHL_BIAS_POWER_SEL = "FALSE",
    parameter PMA_REG_CHL_BIAS_POWER = "FALSE",
    parameter PMA_REG_RX_BUSWIDTH = "40BIT",
    parameter PMA_REG_RX_RATE = "DIV4",
    parameter PMA_REG_RX_RATE_EN = "FALSE",
    parameter integer PMA_REG_RX_RES_TRIM = 55,
    parameter PMA_REG_RX_SIGDET_STATUS_EN = "FALSE",
    parameter integer PMA_REG_CDR_READY_THD_7_0 = 32,
    parameter integer PMA_REG_CDR_READY_THD_11_8 = 0,
    parameter PMA_REG_RX_BUSWIDTH_EN = "FALSE",
    parameter PMA_REG_RX_PCLK_EDGE_SEL = "POS_EDGE",
    parameter integer PMA_REG_CDR_READY_CHECK_CTRL = 0,
    parameter PMA_REG_RX_ICTRL_TRX = "100PCT",
    parameter integer PMA_REG_PRBS_CHK_WIDTH_SEL = 1,
    parameter PMA_REG_RX_ICTRL_PIBUF = "100PCT",
    parameter PMA_REG_RX_ICTRL_PI = "100PCT",
    parameter PMA_REG_RX_ICTRL_DCC = "100PCT",
    parameter PMA_REG_TX_RATE = "DIV1",
    parameter PMA_REG_TX_RATE_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N = "TRUE",
    parameter PMA_REG_RX_TX2RX_PLPBK_RST_N_EN = "FALSE",
    parameter PMA_REG_RX_TX2RX_PLPBK_EN = "FALSE",
    parameter PMA_REG_RX_DATA_POLARITY = "NORMAL",
    parameter PMA_REG_RX_ERR_INSERT = "FALSE",
    parameter PMA_REG_UDP_CHK_EN = "FALSE",
    parameter PMA_REG_PRBS_SEL = "PRBS7",
    parameter PMA_REG_PRBS_CHK_EN = "FALSE",
    parameter integer PMA_REG_LPLL_NFC_STIC_DIS_N = 0,
    parameter PMA_REG_BIST_CHK_PAT_SEL = "PRBS",
    parameter PMA_REG_LOAD_ERR_CNT = "FALSE",
    parameter PMA_REG_CHK_COUNTER_EN = "TRUE",
    parameter integer PMA_REG_CDR_PROP_GAN_SEL = 3,
    parameter integer PMA_REG_CDR_TUBO_PROP_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_GAIN_SEL = 2,
    parameter integer PMA_REG_CDR_TUBO_INT_GAIN_SEL = 6,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_4_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MAX_9_5 = 28,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_2_0 = 0,
    parameter integer PMA_REG_CDR_INT_SAT_MIN_9_3 = 16,
    parameter integer PMA_ANA_RX_REG_O_61_55 = 21,
    parameter integer PMA_ANA_RX_REG_O_69_62 = 0,
    parameter integer PMA_ANA_RX_REG_O_77_70 = 135,
    parameter integer PMA_ANA_RX_REG_O_85_78 = 1,
    parameter integer PMA_ANA_RX_REG_O_93_86 = 8,
    parameter integer PMA_ANA_RX_REG_O_100_94 = 64,
    parameter integer PMA_ANA_RX_REG_O_108_101 = 0,
    parameter integer PMA_ANA_RX_REG_O_111_109 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_4_0 = 3,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MIN_5 = 0,
    parameter integer PMA_REG_OOB_COMWAKE_GAP_MAX = 11,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MIN = 15,
    parameter integer PMA_REG_OOB_COMINIT_GAP_MAX = 35,
    parameter integer PMA_REG_COMWAKE_STATUS_CLEAR = 0,
    parameter integer PMA_REG_COMINIT_STATUS_CLEAR = 0,
    parameter PMA_REG_RX_SATA_COMINIT_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMINIT = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE_OW = "FALSE",
    parameter PMA_REG_RX_SATA_COMWAKE = "FALSE",
    parameter PMA_REG_RX_DCC_DISABLE = "FALSE",
    parameter PMA_REG_RX_SLIP_SEL_EN = "FALSE",
    parameter integer PMA_REG_RX_SLIP_SEL_3_0 = 0,
    parameter PMA_REG_RX_SLIP_EN = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_STATUS_SEL = 5,
    parameter PMA_REG_RX_SIGDET_FSM_RST_N = "TRUE",
    parameter PMA_REG_RX_SIGDET_STATUS = "FALSE",
    parameter PMA_REG_RX_SIGDET_VTH = "36MV",
    parameter integer PMA_REG_RX_SIGDET_GRM = 0,
    parameter PMA_REG_RX_SIGDET_PULSE_EXT = "FALSE",
    parameter integer PMA_REG_RX_SIGDET_CH2_SEL = 0,
    parameter integer PMA_REG_RX_SIGDET_CH2_CHK_WINDOW = 3,
    parameter PMA_REG_RX_SIGDET_CHK_WINDOW_EN = "TRUE",
    parameter integer PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING = 4,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0 = 0,
    parameter integer PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3 = 0,
    parameter integer PMA_REG_RX_SIGDET_4OOB_DET_SEL = 7,
    parameter integer PMA_REG_RX_SIGDET_IC_I = 10,
    parameter integer PMA_REG_RX_EQ1_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ1_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ1_OFF = "FALSE",
    parameter integer PMA_REG_RX_EQ2_R_SET_TOP = 3,
    parameter integer PMA_REG_RX_EQ2_C_SET_FB = 0,
    parameter PMA_REG_RX_EQ2_OFF = "FALSE",
    parameter integer PMA_REG_RX_ICTRL_EQ = 2,
    parameter PMA_REG_EQ_DC_CALIB_EN = "FALSE",
    parameter integer PMA_CTLE_CTRL_REG_I = 0,
    parameter PMA_CTLE_REG_FORCE_SEL_I = "FALSE",
    parameter PMA_CTLE_REG_HOLD_I = "FALSE",
    parameter integer PMA_CTLE_REG_INIT_DAC_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_INIT_DAC_I_3_2 = 0,
    parameter PMA_CTLE_REG_POLARITY_I = "FALSE",
    parameter integer PMA_CTLE_REG_SHIFTER_GAIN_I = 4,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_1_0 = 0,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_9_2 = 1,
    parameter integer PMA_CTLE_REG_THRESHOLD_I_11_10 = 0,
    parameter PMA_REG_RX_RES_TRIM_EN = "FALSE",
    parameter integer PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION = 1,
    parameter integer PMA_REG_ALG_RX_TERM_VCM_SELECTION = 3,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0 = 0,
    parameter integer PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8 = 0,
    parameter PMA_REG_ALG_LOW_SPEED_MODE_ENABLE = "FALSE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER = "TRUE",
    parameter PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION = "FALSE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0 = "TRUE",
    parameter PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1 = "FALSE",
    parameter PMA_REG_EYE_DFETAP1_PLORITY = "FALSE",
    parameter PMA_REG_CDR_SEL = "FALSE",
    parameter PMA_REG_EYE_DET_EN = "FALSE",
    parameter integer PMA_REG_PI_BIAS_CURRENT = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_6_0 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_14_7 = 0,
    parameter integer PMA_REG_ALG_DFE_TEST_SEL_21_15 = 0,
    parameter integer PMA_REG_ALG_EYE_PATH_SEL = 0,
    parameter integer PMA_REG_ALG_CTLE_TEST_SEL = 0,
    parameter PMA_REG_RX_SLIP_SEL_4 = "FALSE",
    parameter PMA_REG_ALG_RX_T1_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_CDRX_BUFF_EN = "TRUE",
    parameter PMA_REG_ALG_RX_VP_T1_SW_PLORITY = "FALSE",
    parameter PMA_REG_ALG_RX_VP_PLORITY = "TRUE",
    parameter PMA_REG_ALG_RX_GAIN_CTRL_SUMMER = "FALSE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_T1_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_VP_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN = "TRUE",
    parameter PMA_REG_ALG_RX_DC_OFFSET_EYE_EN = "TRUE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE = "FALSE",
    parameter PMA_REG_ALG_SLICER_DC_OFFSET_REG = "FALSE",
    parameter PMA_REG_RX_PGA_OFF = "FALSE",
    parameter integer PMA_REG_ALG_CDR_XWEIGHT_I = 4,
    parameter integer PMA_REG_ALG_CDR_YWEIGHT_I = 4,
    parameter PMA_REG_ALG_CTLE_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_CTLE_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_CTLE_INITDAC_6 = 0,
    parameter PMA_REG_ALG_CTLE_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLE_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_2_0 = 4,
    parameter integer PMA_REG_ALG_CTLE_TOPNUM_4_3 = 2,
    parameter PMA_REG_ALG_CTLEOFS_FLIPDIR_I = "TRUE",
    parameter PMA_REG_ALG_CTLEOFS_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_3_0 = 0,
    parameter integer PMA_REG_ALG_CTLEOFS_INITDAC_6_4 = 4,
    parameter PMA_REG_ALG_CTLEOFS_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_CTLEOFS_SHIFT_I = 4,
    parameter PMA_REG_ALG_DFE_CTLE_PWD = "FALSE",
    parameter PMA_REG_ALG_H1_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H1_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_INITDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_H1_INITDAC_6 = 0,
    parameter PMA_REG_ALG_H1_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H1_SHIFT_I = 4,
    parameter PMA_REG_ALG_H2_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H2_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H2_INITDAC_5_1 = 0,
    parameter PMA_REG_ALG_H2_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H2_SHIFT_I_1_0 = 0,
    parameter integer PMA_REG_ALG_H2_SHIFT_I_2 = 1,
    parameter PMA_REG_ALG_H3_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H3_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_INITDAC_4_0 = 0,
    parameter integer PMA_REG_ALG_H3_INITDAC_5 = 1,
    parameter PMA_REG_ALG_H3_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H3_SHIFT_I = 4,
    parameter PMA_REG_ALG_H4_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H4_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_H4_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_H4_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H4_SHIFT_I = 4,
    parameter PMA_REG_ALG_H5_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H5_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_INITDAC = 16,
    parameter PMA_REG_ALG_H5_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H5_SHIFT_I = 4,
    parameter PMA_REG_ALG_H6_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_H6_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_H6_INITDAC_4_3 = 2,
    parameter PMA_REG_ALG_H6_OVERWREN_I = "FALSE",
    parameter integer PMA_REG_ALG_H6_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_HCTLE_OFS_1_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OFS_3_2 = 2,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_5_0 = 0,
    parameter integer PMA_REG_ALG_HCTLE_OVERWRDAC_6 = 1,
    parameter PMA_REG_ALG_HCTLE_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQH_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQH_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQH_REG_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_LEQL_INITDAC_I = 0,
    parameter PMA_REG_ALG_LEQL_PWD_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_REG_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_LEQL_REG_PRESELECT_I = 7,
    parameter integer PMA_REG_ALG_LEQL_REG_SHIFT_I = 4,
    parameter PMA_REG_ALG_NEXTBIT_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_6_0 = 127,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_14_7 = 255,
    parameter integer PMA_REG_ALG_SOFS_COUNTMAX_I_19_15 = 31,
    parameter integer PMA_REG_ALG_SOFS_DACWIN_I = 1,
    parameter PMA_REG_ALG_SOFS_FLIP_DIR_I = "TRUE",
    parameter PMA_REG_ALG_SOFS_FORCE_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_5_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_FORCEDAC_I_6 = 1,
    parameter integer PMA_REG_ALG_SOFS_FORCENUM_I = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_2_0 = 0,
    parameter integer PMA_REG_ALG_SOFS_INITDAC_6_3 = 8,
    parameter integer PMA_REG_ALG_SOFS_SHIFT_I = 1,
    parameter PMA_REG_ALG_SOFS_SKIP_I = "FALSE",
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0 = 254,
    parameter integer PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8 = 15,
    parameter PMA_REG_ALG_ST_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_ST_FORCEN = "FALSE",
    parameter PMA_REG_ALG_ST_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_ST_INITDAC_0 = 0,
    parameter integer PMA_REG_ALG_ST_INITDAC_4_1 = 8,
    parameter PMA_REG_ALG_ST_RECALEN = "FALSE",
    parameter integer PMA_REG_ALG_ST_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_ST_STARTCNT_7_0 = 0,
    parameter integer PMA_REG_ALG_ST_STARTCNT_15_8 = 128,
    parameter integer PMA_REG_ALG_ST_STARTCNT_19_16 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_3_0 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_11_4 = 0,
    parameter integer PMA_REG_ALG_ST_TAPCNT_17_12 = 2,
    parameter integer PMA_REG_ALG_ST_TOPTAP_1_0 = 3,
    parameter integer PMA_REG_ALG_ST_TOPTAP_3_2 = 3,
    parameter integer PMA_REG_ALG_SWCLK_DIV = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_3_0 = 0,
    parameter integer PMA_REG_ALG_TAPA_DAC_4 = 1,
    parameter integer PMA_REG_ALG_TAPA_NUM = 7,
    parameter integer PMA_REG_ALG_TAPB_DAC_0 = 0,
    parameter integer PMA_REG_ALG_TAPB_DAC_4_1 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_3_0 = 8,
    parameter integer PMA_REG_ALG_TAPB_NUM_5_4 = 0,
    parameter integer PMA_REG_ALG_TAPC_DAC = 16,
    parameter integer PMA_REG_ALG_TAPC_NUM_0 = 1,
    parameter integer PMA_REG_ALG_TAPC_NUM_5_1 = 4,
    parameter integer PMA_REG_ALG_TAPD_DAC_2_0 = 0,
    parameter integer PMA_REG_ALG_TAPD_DAC_4_3 = 2,
    parameter integer PMA_REG_ALG_TAPD_NUM = 10,
    parameter PMA_REG_ALG_VP_FLIPDIR_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_GRN_SHIFT_I = 5,
    parameter PMA_REG_ALG_VP_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_VP_IDEAL_2_0 = 0,
    parameter integer PMA_REG_ALG_VP_IDEAL_6_3 = 10,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_3_0 = 0,
    parameter integer PMA_REG_ALG_VP_INITDAC_I_6_4 = 0,
    parameter PMA_REG_ALG_VP_OVERWREN = "FALSE",
    parameter integer PMA_REG_ALG_VP_RED_SHIFT_I = 5,
    parameter integer PMA_REG_ALG_VPOFS_SEL_0 = 0,
    parameter integer PMA_REG_ALG_VPOFS_SEL_2_1 = 1,
    parameter integer PMA_REG_ALG_H1_UPBOUND_5_0 = 55,
    parameter integer PMA_REG_ALG_H1_UPBOUND_6 = 1,
    parameter PMA_REG_ALG_CTLEOFS_PWDN = "FALSE",
    parameter PMA_REG_ALG_LEQH_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_LEQL_OVEREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_FLIPDIR_I = "FALSE",
    parameter PMA_REG_ALG_AGC_HOLD_I = "FALSE",
    parameter integer PMA_REG_ALG_AGC_INITDAC = 10,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_1_0 = 3,
    parameter integer PMA_REG_ALG_AGC_LOWBOUND_3_2 = 0,
    parameter PMA_REG_ALG_AGC_OVERWREN_I = "FALSE",
    parameter PMA_REG_ALG_AGC_PWD = "FALSE",
    parameter integer PMA_REG_ALG_AGC_SHIFT_I = 4,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_0 = 1,
    parameter integer PMA_REG_ALG_AGC_UPBOUND_3_1 = 7,
    parameter integer PMA_REG_ALG_AGC_WAITSEL = 11,
    parameter PMA_REG_PI_CTRL_SEL_RX = "FALSE",
    parameter integer PMA_REG_PI_CTRL_RX_4_0 = 0,
    parameter integer PMA_REG_PI_CTRL_RX_7_5 = 0,
    parameter PMA_CFG_RX_LANE_POWERUP = "ON",
    parameter PMA_CFG_RX_PMA_RSTN = "TRUE",
    parameter PMA_INT_PMA_RX_MASK_0 = "FALSE",
    parameter PMA_INT_PMA_RX_CLR_0 = "FALSE",
    parameter PMA_CFG_CTLE_ADP_RSTN = "TRUE",
    parameter PMA_CFG_RX_CDR_RSTN = "TRUE",
    parameter PMA_CFG_RX_CLKPATH_RSTN = "TRUE",
    parameter PMA_CFG_RX_DFE_RSTN = "TRUE",
    parameter PMA_CFG_RX_LEQ_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIDING_RSTN = "TRUE",
    parameter PMA_CFG_RX_EYE_RSTN = "TRUE",
    parameter PMA_CFG_RX_CTLE_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLICER_DCCAL_RSTN = "TRUE",
    parameter PMA_CFG_RX_SLIP_RSTN = "TRUE",
    parameter integer PMA_REG_TX_BEACON_TIMER_SEL = 0,
    parameter PMA_REG_TX_BIT_CONV = "FALSE",
    parameter integer PMA_REG_TX_RES_CAL = 50,
    parameter integer PMA_REG_TX_UDP_DATA_20 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_26_21 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_34_27 = 0,
    parameter integer PMA_REG_TX_UDP_DATA_39_25 = 0,
    parameter integer PMA_REG_TX_BUSWIDTH_EN = 0,
    parameter PMA_REG_TX_PD_POST = "OFF",
    parameter PMA_REG_TX_PD_POST_OW = "FALSE",
    parameter PMA_REG_TX_BUSWIDTH = "20BIT",
    parameter integer PMA_REG_EI_PCLK_DELAY_SEL = 0,
    parameter integer PMA_REG_TX_AMP_DAC0 = 25,
    parameter integer PMA_REG_TX_AMP_DAC1 = 19,
    parameter integer PMA_REG_TX_AMP_DAC2 = 14,
    parameter integer PMA_REG_TX_AMP_DAC3 = 9,
    parameter PMA_REG_TX_RXDET_THRESHOLD = "84MV",
    parameter PMA_REG_TX_BEACON_OSC_CTRL = "FALSE",
    parameter integer PMA_REG_TX_PRBS_GEN_WIDTH_SEL = 0,
    parameter PMA_REG_TX_TX2RX_SLPBACK_EN = "FALSE",
    parameter PMA_REG_TX_PCLK_EDGE_SEL = "FALSE",
    parameter PMA_REG_TX_PRBS_GEN_EN = "FALSE",
    parameter PMA_REG_TX_PRBS_SEL = "PRBS7",
    parameter integer PMA_REG_TX_UDP_DATA_7_TO_0 = 5,
    parameter integer PMA_REG_TX_UDP_DATA_15_TO_8 = 235,
    parameter integer PMA_REG_TX_UDP_DATA_19_TO_16 = 3,
    parameter integer PMA_REG_TX_FIFO_WP_CTRL = 4,
    parameter PMA_REG_TX_FIFO_EN = "FALSE",
    parameter integer PMA_REG_TX_DATA_MUX_SEL = 0,
    parameter PMA_REG_TX_ERR_INSERT = "FALSE",
    parameter PMA_REG_TX_SATA_EN = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON_OW = "FALSE",
    parameter PMA_REG_RATE_CHANGE_TXPCLK_ON = "TRUE",
    parameter integer PMA_REG_TX_CFG_POST1 = 0,
    parameter integer PMA_REG_TX_CFG_POST2 = 0,
    parameter integer PMA_REG_TX_OOB_DELAY_SEL = 0,
    parameter PMA_REG_TX_POLARITY = "NORMAL",
    parameter PMA_REG_TX_LS_MODE_EN = "FALSE",
    parameter PMA_REG_RX_JTAG_OE = "TRUE",
    parameter integer PMA_REG_RX_ACJTAG_VHYSTSEL = 0,
    parameter PMA_REG_TX_RES_CAL_EN = "FALSE",
    parameter integer PMA_REG_RX_TERM_MODE_CTRL = 5,
    parameter PMA_REG_PLPBK_TXPCLK_EN = "FALSE",
    parameter integer PMA_REG_TX_PH_SEL_0 = 1,
    parameter integer PMA_REG_TX_PH_SEL_6_1 = 0,
    parameter integer PMA_REG_TX_CFG_PRE = 0,
    parameter integer PMA_REG_TX_CFG_MAIN = 0,
    parameter integer PMA_REG_CFG_POST = 0,
    parameter PMA_REG_PD_MAIN = "TRUE",
    parameter PMA_REG_PD_PRE = "TRUE",
    parameter integer PMA_REG_TX_RXDET_TIMER_SEL = 87,
    parameter PMA_REG_TX_MOD_STAND_BY_EN = "FALSE",
    parameter PMA_REG_STATE_STAND_BY_SEL = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW = "FALSE",
    parameter PMA_REG_TX_SYNC_NEW_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_OW = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_POLAR_CTRL = "FALSE",
    parameter PMA_REG_TX_FREERUN_PD = "TRUE",
    parameter PMA_REG_TX_CHANGE_ON_SEL = "FALSE",
    parameter PMA_REG_TX_CHANGE_ON_CTRL = "FALSE",
    parameter integer PMA_REG_TX_FREERUN_RATE_0 = 0,
    parameter integer PMA_REG_TX_FREERUN_RATE_1 = 0,
    parameter PMA_REG_TX_FREERUN_RATE_OW = "FALSE",
    parameter PMA_REG_TX_RST_SYNC_CLK_SEL = "TRUE",
    parameter integer PMA_REG_TX_PI_CTRL_SEL = 0,
    parameter integer PMA_REG_TX_PI_CTRL = 0,
    parameter PMA_LANE_POWERUP = "TRUE",
    parameter PMA_POR_N = "TRUE",
    parameter PMA_TX_LANE_POWERUP = "TRUE",
    parameter PMA_TX_PMA_RSTN = "TRUE",
    parameter PMA_LPLL_POWERUP = "TRUE",
    parameter PMA_LPLL_RSTN = "TRUE",
    parameter PMA_LPLL_LOCKDET_RSTN = "TRUE",
    parameter integer PMA_REG_LPLL_PFDDELAY_SEL = 1,
    parameter PMA_REG_LPLL_PFDDELAY_EN = "TRUE",
    parameter integer PMA_REG_LPLL_VCTRL_SET = 0,
    parameter PMA_LPLL_CHARGE_PUMP_CTRL = "type",
    parameter PMA_LPLL_REFDIV = "DIV1",
    parameter integer PMA_LPLL_FBDIV = 38,
    parameter integer PMA_LPLL_LPF_RES = 1,
    parameter integer PMA_LPLL_REFLOSS_READY = 0,
    parameter integer PMA_LPLL_LOCKED_PFDDELAY = 0,
    parameter integer PMA_LPLL_MCLK_SEL = 0,
    parameter integer PMA_LPLL_TEST_SEL = 0,
    parameter PMA_LPLL_TEST_SIG_HALF_EN = "TRUE",
    parameter PMA_LPLL_TEST_V_EN = "FALSE",
    parameter PMA_LPLL_MCLK_EN = "TRUE",
    parameter integer PMA_LPLL_MCLK_DET_CTL = 16,
    parameter integer PMA_LPLL_LOCKDET_REFCT = 3,
    parameter integer PMA_LPLL_LOCKDET_FBCT = 3,
    parameter integer PMA_LPLL_LOCKDET_LOCKCT = 4,
    parameter integer PMA_LPLL_LOCKDET_ITER = 1,
    parameter integer PMA_LPLL_UNLOCKDET_ITER = 2,
    parameter integer PMA_LPLL_LOCKDET_EN_OW = 0,
    parameter integer PMA_LPLL_LOCKDET_EN = 0,
    parameter integer PMA_LPLL_LOCKDET_MODE = 0,
    parameter integer PMA_LPLL_LOCKDET_OW = 0,
    parameter integer PMA_LPLL_LOCKDETED = 0,
    parameter integer PMA_LPLL_UNLOCKDET_OW = 0,
    parameter integer PMA_LPLL_UNLOCKDETED = 0,
    parameter integer PMA_LPLL_LOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_UNLOCKED_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_LOCKDET_REPEAT = 0,
    parameter integer PMA_LPLL_NOFBCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_NOREFCLK_STICKY_CLEAR = 0,
    parameter integer PMA_LPLL_READY_OR_LOCK = 0,
    parameter integer PMA_LPLL_READY = 0,
    parameter integer PMA_LPLL_READY_OW = 0,
    parameter PMA_REG_TXCLK_SEL = "HPLL",
    parameter PMA_REG_RXCLK_SEL = "HPLL",
    parameter integer PMA_REG_TEST_BUF = 0,
    parameter integer PMA_REG_CHL_TEST = 0
) (
    output P_CFG_READY,
    output [7:0] P_CFG_RDATA,
    output P_CFG_INT,
    output [24:0] LANE_COUT_BUS_FORWARD,
    output [1:0] LANE_COUT_BUS_BACKWARD,
    output P_RX_PRBS_ERROR,
    output P_PCS_RX_MCB_STATUS,
    output P_PCS_LSM_SYNCED,
    output [87:0] P_RDATA,
    output P_RXDVLD,
    output P_RXDVLD_H,
    output [5:0] P_RXSTATUS,
    output [2:0] P_EM_ERROR_CNT,
    output P_LPLL_READY,
    output P_RX_SIGDET_STATUS,
    output P_RX_SATA_COMINIT,
    output P_RX_SATA_COMWAKE,
    output P_RX_LS_DATA,
    output P_RX_READY,
    output [19:0] P_TEST_STATUS,
    output P_TX_RXDET_STATUS,
    output P_RCLK2FABRIC,
    output P_TCLK2FABRIC,
    output P_CA_ALIGN_RX,
    output P_CA_ALIGN_TX,
    output P_TX_SDN,
    output P_TX_SDP,
    input P_RX_CLK_FR_CORE,
    input P_RCLK2_FR_CORE,
    input P_TX_CLK_FR_CORE,
    input P_TCLK2_FR_CORE,
    input P_PCS_RX_RST,
    input P_PCS_TX_RST,
    input P_EXT_BRIDGE_PCS_RST,
    input P_CFG_RST,
    input P_CFG_CLK,
    input P_CFG_PSEL,
    input P_CFG_ENABLE,
    input P_CFG_WRITE,
    input [11:0] P_CFG_ADDR,
    input [7:0] P_CFG_WDATA,
    input [24:0] LANE_CIN_BUS_FORWARD,
    input [1:0] LANE_CIN_BUS_BACKWARD,
    input [87:0] P_TDATA,
    input P_PCIE_EI_H,
    input P_PCIE_EI_L,
    input [15:0] P_TX_DEEMP,
    input [1:0] P_TX_DEEMP_POST_SEL,
    input P_BLK_ALIGN_CTRL,
    input P_TX_ENC_TYPE,
    input P_RX_DEC_TYPE,
    input P_PCS_BIT_SLIP,
    input P_PCS_WORD_ALIGN_EN,
    input P_RX_POLARITY_INVERT,
    input P_PCS_MCB_EXT_EN,
    input P_PCS_NEAREND_LOOP,
    input P_PCS_FAREND_LOOP,
    input P_PMA_NEAREND_PLOOP,
    input P_PMA_NEAREND_SLOOP,
    input P_PMA_FAREND_PLOOP,
    input P_PCS_PRBS_EN,
    input P_LANE_POWERDOWN,
    input P_LANE_RST,
    input P_RX_LANE_POWERDOWN,
    input P_RX_PMA_RST,
    input P_RX_CDR_RST,
    input P_RX_CLKPATH_RST,
    input P_RX_DFE_RST,
    input P_RX_LEQ_RST,
    input P_RX_SLIDING_RST,
    input P_RX_DFE_EN,
    input P_RX_T1_EN,
    input P_RX_CDRX_EN,
    input P_RX_T1_DFE_EN,
    input P_RX_T2_DFE_EN,
    input P_RX_T3_DFE_EN,
    input P_RX_T4_DFE_EN,
    input P_RX_T5_DFE_EN,
    input P_RX_T6_DFE_EN,
    input P_RX_SLIDING_EN,
    input P_RX_EYE_RST,
    input P_RX_EYE_EN,
    input [7:0] P_RX_EYE_TAP,
    input [7:0] P_RX_PIC_EYE,
    input [7:0] P_RX_PIC_FASTLOCK,
    input P_RX_PIC_FASTLOCK_STROBE,
    input P_EM_RD_TRIGGER,
    input [1:0] P_EM_MODE_CTRL,
    input P_RX_CTLE_DCCAL_RST,
    input P_RX_SLICER_DCCAL_RST,
    input P_RX_SLICER_DCCAL_EN,
    input P_RX_CTLE_DCCAL_EN,
    input P_RX_SLIP_RST,
    input P_RX_SLIP_EN,
    input P_LPLL_POWERDOWN,
    input P_LPLL_RST,
    input P_LPLL_LOCKDET_RST,
    input P_TX_LS_DATA,
    input P_TX_BEACON_EN,
    input P_TX_SWING,
    input P_TX_RXDET_REQ,
    input [1:0] P_TX_RATE,
    input [2:0] P_TX_BUSWIDTH,
    input [2:0] P_TX_FREERUN_BUSWIDTH,
    input [2:0] P_TX_MARGIN,
    input P_TX_PMA_RST,
    input P_TX_LANE_POWERDOWN,
    input P_TX_PIC_EN,
    input [1:0] P_RX_RATE,
    input [2:0] P_RX_BUSWIDTH,
    input P_RX_HIGHZ,
    input [7:0] P_CIM_CLK_ALIGNER_RX,
    input [7:0] P_CIM_CLK_ALIGNER_TX,
    input P_ALIGN_MODE_VALID_RX,
    input [1:0] P_ALIGN_MODE_RX,
    input P_ALIGN_MODE_VALID_TX,
    input [2:0] P_ALIGN_MODE_TX,
    input PMA_HPLL_CK0,
    input PMA_HPLL_CK90,
    input PMA_HPLL_CK180,
    input PMA_HPLL_CK270,
    input PMA_HPLL_READY_IN,
    input PMA_HPLL_REFCLK_IN,
    input [1:0] PMA_IPN50U_IN,
    input PMA_LPLL_REFCLK,
    input [5:0] PMA_RES_CAL_I,
    input PMA_TX_SYNC_HPLL,
    input PMA_TX_RATE_CHANGE_ON_0,
    input PMA_TX_RATE_CHANGE_ON_1,
    input PMA_TX_SYNC,
    input P_RX_SDN,
    input P_RX_SDP
)  ;
endmodule


module GTP_IDDR_E1
#(
    parameter GRS_EN = "TRUE",
    parameter IDDR_MODE = "OPPOSITE_EDGE",
    parameter RS_TYPE = "ASYNC_RESET"
) (
    output Q0,
    output Q1,
    input D,
    input CLK,
    input CE,
    input RS
)  ;
endmodule


module GTP_INBUF
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    input I
)  ;
endmodule


module GTP_INBUFDS
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    input I,
    input IB
)  ;
endmodule


module GTP_INBUFDS_E1
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    output OB,
    input I,
    input IB
)  ;
endmodule


module GTP_INBUFE
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    input EN,
    input I
)  ;
endmodule


module GTP_INBUFEDS
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    input EN,
    input I,
    input IB
)  ;
endmodule


module GTP_INBUFEDS_E1
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    output OB,
    input EN,
    input I,
    input IB
)  ;
endmodule


module GTP_INBUFG
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    input I
)  ;
endmodule


module GTP_INBUFGDS
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    input I,
    input IB
)  ;
endmodule


module GTP_INV
(
    output Z,
    input I
)  ;
endmodule


module GTP_IOBUF
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8",
    parameter TERM_DDR = "ON"
) (
    output O,
    inout IO,
    input I,
    input T
)  ;
endmodule


module GTP_IOBUF_RX_MIPI
#(
    parameter HPIO = "FALSE",
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "6",
    parameter TERM_DIFF = "ON"
) (
    output O_LP,
    output OB_LP,
    output O_HS,
    inout IO,
    inout IOB,
    input I_LP,
    input IB_LP,
    input T,
    input TB,
    input M
)  ;
endmodule


module GTP_IOBUF_TX_MIPI
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "6",
    parameter TERM_DIFF = "ON"
) (
    output O_LP,
    output OB_LP,
    inout IO,
    inout IOB,
    input I_LP,
    input IB_LP,
    input I_HS,
    input T,
    input TB,
    input M
)  ;
endmodule


module GTP_IOBUFCO
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    inout IO,
    inout IOB,
    input I,
    input T
)  ;
endmodule


module GTP_IOBUFCO_E1
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    inout IO,
    inout IOB,
    input I,
    input IB,
    input T,
    input TB
)  ;
endmodule


module GTP_IOBUFDS
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    inout IO,
    inout IOB,
    input I,
    input T
)  ;
endmodule


module GTP_IOBUFE
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8",
    parameter TERM_DDR = "ON"
) (
    output O,
    inout IO,
    input I,
    input EN,
    input T
)  ;
endmodule


module GTP_IOBUFECO
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DDR = "ON"
) (
    output O,
    inout IO,
    inout IOB,
    input I,
    input EN,
    input T
)  ;
endmodule


module GTP_IOBUFEDS
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter TERM_DIFF = "ON"
) (
    output O,
    inout IO,
    inout IOB,
    input I,
    input EN,
    input T
)  ;
endmodule


module GTP_IOCLKBUF
#(
    parameter GATE_EN = "FALSE"
) (
    output CLKOUT,
    input CLKIN,
    input DI
)  ;
endmodule


module GTP_IOCLKDIV_E2
#(
    parameter DIV_FACTOR = "BYPASS"
) (
    output CLKDIVOUT,
    input CLKIN,
    input RST_N,
    input CE
)  ;
endmodule


module GTP_IOCLKDIV_E3
#(
    parameter DIV_FACTOR = "8",
    parameter PHASE_SHIFT = "0"
) (
    input RST,
    input CLKIN,
    output CLKDIVOUT
)  ;
endmodule


module GTP_IODELAY_E2
#(
    parameter [7:0] DELAY_STEP_VALUE = 8'h00,
    parameter DELAY_STEP_SEL = "PARAMETER",
    parameter TDELAY_EN = "FALSE"
) (
    output DO,
    input DI,
    input DELAY_SEL,
    input [7:0] DELAY_STEP,
    input EN_N
)  ;
endmodule


module GTP_IPAL_E2
#(
    parameter DATA_WIDTH = "X8",
    parameter [31:0] IDCODE = 32'hAAAA5555,
    parameter SIM_DEVICE = "PG2L100H"
) (
    output [31:0] DO,
    output RBCRC_ERR,
    output RBCRC_VALID,
    output ECC_VALID,
    output [11:0] ECC_INDEX,
    output SERROR,
    output DERROR,
    output [7:0] SEU_FRAME_ADDR,
    output [7:0] SEU_COLUMN_ADDR,
    output [4:0] SEU_REGION_ADDR,
    output [7:0] SEU_FRAME_NADDR,
    output [7:0] SEU_COLUMN_NADDR,
    output [4:0] SEU_REGION_NADDR,
    output PRCFG_OVER,
    output PRCFG_ERR,
    output DRCFG_OVER,
    output DRCFG_ERR,
    input RST_N,
    input CLK,
    input CS_N,
    input RW_SEL,
    input [31:0] DI
)  ;
endmodule


module GTP_ISERDES_E2
#(
    parameter ISERDES_MODE = "SDR1TO4",
    parameter GRS_EN = "TRUE",
    parameter CASCADE_MODE = "MASTER",
    parameter BITSLIP_EN = "FALSE",
    parameter integer NUM_ICE = 0,
    parameter GRS_TYPE_Q0 = "RESET",
    parameter GRS_TYPE_Q1 = "RESET",
    parameter GRS_TYPE_Q2 = "RESET",
    parameter GRS_TYPE_Q3 = "RESET",
    parameter LRS_TYPE_Q0 = "ASYNC_RESET",
    parameter LRS_TYPE_Q1 = "ASYNC_RESET",
    parameter LRS_TYPE_Q2 = "ASYNC_RESET",
    parameter LRS_TYPE_Q3 = "ASYNC_RESET",
    parameter HPIO = "FALSE"
) (
    input RST,
    input ICE0,
    input ICE1,
    input DESCLK,
    input ICLK,
    input ICLKB,
    input OCLK,
    input ICLKDIV,
    input DI,
    input BITSLIP,
    input ISHIFTIN0,
    input ISHIFTIN1,
    input [2:0] IFIFO_WADDR,
    input [2:0] IFIFO_RADDR,
    output [7:0] DO,
    output ISHIFTOUT0,
    output ISHIFTOUT1
)  ;
endmodule


module GTP_ISERDES_FIFO
#(
    parameter FIFO_BYPASS = "FALSE",
    parameter WCLK_INV = "FALSE",
    parameter RCLK_INV = "FALSE"
) (
    output [7:0] DOUT,
    output VALID_O,
    input [7:0] DIN,
    input VALID_I,
    input RST,
    input EN,
    input WCLK,
    input RCLK,
    output EMPTY,
    output FULL
)  ;
endmodule


module GTP_JTAGIF
#(
    parameter [31:0] USERCODE = 32'hFFFFFFFF,
    parameter [31:0] IDCODE = 32'h5555AAAA
) (
    output TDO,
    input TCK,
    input TMS,
    input TDI
)  ;
endmodule


module GTP_KEYRAM
(
    input ERASE_KEY_N
)  ;
endmodule


module GTP_LUT1
#(
    parameter [1:0] INIT = 2'h0
) (
    output Z,
    input I0
)  ;
endmodule


module GTP_LUT2
#(
    parameter [3:0] INIT = 4'h0
) (
    output Z,
    input I0,
    input I1
)  ;
endmodule


module GTP_LUT3
#(
    parameter [7:0] INIT = 8'h00
) (
    output Z,
    input I0,
    input I1,
    input I2
)  ;
endmodule


module GTP_LUT4
#(
    parameter [15:0] INIT = 16'h0000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3
)  ;
endmodule


module GTP_LUT5
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4
)  ;
endmodule


module GTP_LUT6
#(
    parameter [63:0] INIT = 64'h0000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5
)  ;
endmodule


module GTP_LUT6CARRY
#(
    parameter [63:0] INIT = 64'h0000000000000000,
    parameter I5_TO_CARRY = "TRUE",
    parameter I5_TO_LUT = "FALSE"
) (
    output COUT,
    output Z,
    input CIN,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5
)  ;
endmodule


module GTP_LUT6D
#(
    parameter [63:0] INIT = 64'h0000000000000000
) (
    output Z,
    output Z5,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5
)  ;
endmodule


module GTP_LUT7
#(
    parameter [127:0] INIT = 128'h00000000000000000000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5,
    input I6
)  ;
endmodule


module GTP_LUT8
#(
    parameter [255:0] INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5,
    input I6,
    input I7
)  ;
endmodule


module GTP_MONITOR_E1
#(
    parameter MODE = "DEFAULT",
    parameter CALIB = "FALSE",
    parameter DYN_CALIB = "FALSE",
    parameter integer AVG_NUM = 16,
    parameter [1:0] SAMPLE_AL = 2'h0
) (
    input RST_N,
    input CLK,
    input EN,
    input SAMPLE,
    input [4:0] SEL,
    output [9:0] DATA,
    output DATA_VALID,
    output READY
)  ;
endmodule


module GTP_MONITOR_E1_DFT
#(
    parameter [11:0] ANA_INIT = 12'h00f,
    parameter [4:0] DATA_COUNT = 5'h0d,
    parameter MODE = "DEFAULT",
    parameter CALIB = "FALSE",
    parameter DYN_CALIB = "FALSE",
    parameter integer AVG_NUM = 16,
    parameter TEST_JTAG_EN = "FALSE",
    parameter [1:0] SAMPLE_AL = 2'h0
) (
    input RST_N,
    input CLK,
    input EN,
    input SAMPLE,
    input [4:0] SEL,
    input TEST_BIST_MODE,
    input TEST_BIST_START,
    input TEST_TDI,
    input TEST_TCK,
    input TEST_FLG_JTAG,
    input TEST_SHIFTDR,
    input TEST_CLOCKDR,
    input TEST_CAPTUREDR,
    input TEST_UPDATEDR,
    input [9:0] TEST_BIST_REF_MAX,
    input [9:0] TEST_BIST_REF_MIN,
    output [9:0] DATA,
    output DATA_VALID,
    output READY,
    output TEST_TDO,
    output TEST_BIST_VALID,
    output TEST_BIST_ERROR
)  ;
endmodule


module GTP_MUX2LUT7
(
    output Z,
    input I0,
    input I1,
    input S
)  ;
endmodule


module GTP_MUX2LUT8
(
    output Z,
    input I0,
    input I1,
    input S
)  ;
endmodule


module GTP_ODDR_E1
#(
    parameter GRS_EN = "TRUE",
    parameter ODDR_MODE = "SAME_EDGE",
    parameter RS_TYPE = "ASYNC_RESET"
) (
    output Q,
    input D0,
    input D1,
    input CLK,
    input CE,
    input RS
)  ;
endmodule


module GTP_ONE
(
    output Z
)  ;
endmodule


module GTP_OSC_E4
(
    output CLKOUT,
    input EN_N
)  ;
endmodule


module GTP_OSERDES_E2
#(
    parameter GRS_EN = "TRUE",
    parameter OSERDES_MODE = "SDR4TO1",
    parameter TSERDES_EN = "FALSE",
    parameter UPD0_SHIFT_EN = "FALSE",
    parameter UPD1_SHIFT_EN = "FALSE",
    parameter [1:0] INIT_SET = 2'b00,
    parameter GRS_TYPE_DQ = "RESET",
    parameter LRS_TYPE_DQ0 = "ASYNC_RESET",
    parameter LRS_TYPE_DQ1 = "ASYNC_RESET",
    parameter LRS_TYPE_DQ2 = "ASYNC_RESET",
    parameter LRS_TYPE_DQ3 = "ASYNC_RESET",
    parameter GRS_TYPE_TQ = "RESET",
    parameter LRS_TYPE_TQ0 = "ASYNC_RESET",
    parameter LRS_TYPE_TQ1 = "ASYNC_RESET",
    parameter LRS_TYPE_TQ2 = "ASYNC_RESET",
    parameter LRS_TYPE_TQ3 = "ASYNC_RESET",
    parameter TRI_EN = "FALSE",
    parameter TBYTE_EN = "FALSE",
    parameter MIPI_EN = "FALSE",
    parameter OCASCADE_EN = "FALSE",
    parameter HPIO = "FALSE",
    parameter ODELAY_EN = "FALSE",
    parameter TDELAY_EN = "FALSE",
    parameter TSERDES_MODE = "SDR4TO1",
    parameter TUPD0_SHIFT_EN = "FALSE",
    parameter TUPD1_SHIFT_EN = "FALSE",
    parameter [1:0] TINIT_SET = 2'b00,
    parameter TERMBYTE_EN = "FALSE",
    parameter TERM_EN = "FALSE",
    parameter [1:0] TERM_OFF_SET = 2'b00,
    parameter [1:0] TERM_ON_SET = 2'b00
) (
    input RST,
    input OCE,
    input TCE,
    input OCLKDIV,
    input SERCLK,
    input OCLK,
    input MIPI_CTRL,
    input UPD0_SHIFT,
    input UPD1_SHIFT,
    input OSHIFTIN0,
    input OSHIFTIN1,
    input [7:0] DI,
    input [7:0] TI,
    input TBYTE_IN,
    output OSHIFTOUT0,
    output OSHIFTOUT1,
    output TQ,
    output DO,
    output TFB,
    output TERM_FB
)  ;
endmodule


module GTP_OSERDES_FIFO
#(
    parameter FIFO_BYPASS = "FASLE",
    parameter WCLK_INV = "FALSE",
    parameter RCLK_INV = "FALSE"
) (
    output [7:0] DOUT,
    output [7:0] TOUT,
    input [7:0] DIN,
    input [7:0] TIN,
    input RST,
    input EN,
    input WCLK,
    input RCLK,
    output EMPTY,
    output FULL
)  ;
endmodule


module GTP_OUTBUF
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8"
) (
    output O,
    input I
)  ;
endmodule


module GTP_OUTBUFCO
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I
)  ;
endmodule


module GTP_OUTBUFCO_E1
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I,
    input IB
)  ;
endmodule


module GTP_OUTBUFDS
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I
)  ;
endmodule


module GTP_OUTBUFT
#(
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW_RATE = "SLOW",
    parameter DRIVE_STRENGTH = "8"
) (
    output O,
    input I,
    input T
)  ;
endmodule


module GTP_OUTBUFTCO
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I,
    input T
)  ;
endmodule


module GTP_OUTBUFTCO_E1
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I,
    input IB,
    input T,
    input TB
)  ;
endmodule


module GTP_OUTBUFTDS
#(
    parameter IOSTANDARD = "DEFAULT"
) (
    output O,
    output OB,
    input I,
    input T
)  ;
endmodule


module GTP_PCIEGEN2
#(
    parameter GRS_EN = "TRUE",
    parameter PIN_MUX_INT_FORCE_EN = "FALSE",
    parameter PIN_MUX_INT_DISABLE = "FALSE",
    parameter DIAG_CTRL_BUS_B2 = "NORMAL",
    parameter DYN_DEBUG_SEL_EN = "FALSE",
    parameter integer DEBUG_INFO_SEL = 0,
    parameter integer BAR_RESIZABLE = 21,
    parameter integer NUM_OF_RBARS = 3,
    parameter integer BAR_INDEX_0 = 0,
    parameter integer BAR_INDEX_1 = 2,
    parameter integer BAR_INDEX_2 = 4,
    parameter TPH_DISABLE = "FALSE",
    parameter MSIX_CAP_DISABLE = "FALSE",
    parameter MSI_CAP_DISABLE = "FALSE",
    parameter MSI_PVM_DISABLE = "FALSE",
    parameter integer BAR_MASK_WRITABLE = 32,
    parameter integer APP_DEV_NUM = 0,
    parameter integer APP_BUS_NUM = 0,
    parameter RAM_MUX_EN = "FALSE",
    parameter ATOMIC_DISABLE = "FALSE"
) (
    input MEM_CLK,
    input PCLK,
    input PCLK_DIV2,
    input BUTTON_RST,
    input POWER_UP_RST,
    input PERST,
    output CORE_RST_N,
    output TRAINING_RST_N,
    input APP_INIT_RST,
    output PHY_RST_N,
    input [2:0] DEVICE_TYPE,
    input RX_LANE_FLIP_EN,
    input TX_LANE_FLIP_EN,
    input APP_LTSSM_EN,
    output SMLH_LINK_UP,
    output RDLH_LINK_UP,
    input APP_REQ_RETRY_EN,
    output [4:0] SMLH_LTSSM_STATE,
    output AXIS_MASTER_TVALID,
    input AXIS_MASTER_TREADY,
    output [127:0] AXIS_MASTER_TDATA,
    output [3:0] AXIS_MASTER_TKEEP,
    output AXIS_MASTER_TLAST,
    output [7:0] AXIS_MASTER_TUSER,
    input [2:0] TRGT1_RADM_PKT_HALT,
    output [5:0] RADM_GRANT_TLP_TYPE,
    output AXIS_SLAVE0_TREADY,
    input AXIS_SLAVE0_TVALID,
    input [127:0] AXIS_SLAVE0_TDATA,
    input AXIS_SLAVE0_TLAST,
    input AXIS_SLAVE0_TUSER,
    output AXIS_SLAVE1_TREADY,
    input AXIS_SLAVE1_TVALID,
    input [127:0] AXIS_SLAVE1_TDATA,
    input AXIS_SLAVE1_TLAST,
    input AXIS_SLAVE1_TUSER,
    output AXIS_SLAVE2_TREADY,
    input AXIS_SLAVE2_TVALID,
    input [127:0] AXIS_SLAVE2_TDATA,
    input AXIS_SLAVE2_TLAST,
    input AXIS_SLAVE2_TUSER,
    output PM_XTLH_BLOCK_TLP,
    input [31:0] DBI_ADDR,
    input [31:0] DBI_DIN,
    input DBI_CS,
    input DBI_CS2,
    input [3:0] DBI_WR,
    input APP_DBI_RO_WR_DISABLE,
    output LBC_DBI_ACK,
    output [31:0] LBC_DBI_DOUT,
    output SEDO,
    output SEDO_EN,
    input SEDI,
    input SEDI_ACK,
    output CFG_INT_DISABLE,
    input SYS_INT,
    output INTA_GRT_MUX,
    output INTB_GRT_MUX,
    output INTC_GRT_MUX,
    output INTD_GRT_MUX,
    input VEN_MSI_REQ,
    input [2:0] VEN_MSI_TC,
    input [4:0] VEN_MSI_VECTOR,
    output VEN_MSI_GRANT,
    input [31:0] CFG_MSI_PENDING,
    output CFG_MSI_EN,
    input [63:0] MSIX_ADDR,
    input [31:0] MSIX_DATA,
    output CFG_MSIX_EN,
    output CFG_MSIX_FUNC_MASK,
    output RADM_PM_TURNOFF,
    output RADM_MSG_UNLOCK,
    input OUTBAND_PWRUP_CMD,
    output PM_STATUS,
    output [2:0] PM_DSTATE,
    output AUX_PM_EN,
    output PM_PME_EN,
    output PM_LINKST_IN_L0S,
    output PM_LINKST_IN_L1,
    output PM_LINKST_IN_L2,
    output PM_LINKST_L2_EXIT,
    input APP_REQ_ENTR_L1,
    input APP_READY_ENTR_L23,
    input APP_REQ_EXIT_L1,
    input APP_XFER_PENDING,
    output WAKE,
    output RADM_PM_PME,
    output RADM_PM_TO_ACK,
    input APPS_PM_XMT_TURNOFF,
    input APP_UNLOCK_MSG,
    input APPS_PM_XMT_PME,
    input APP_CLK_PM_EN,
    output [4:0] PM_MASTER_STATE,
    output [4:0] PM_SLAVE_STATE,
    input SYS_AUX_PWR_DET,
    input APP_HDR_VALID,
    input [127:0] APP_HDR_LOG,
    input [12:0] APP_ERR_BUS,
    input APP_ERR_ADVISORY,
    output CFG_SEND_COR_ERR_MUX,
    output CFG_SEND_NF_ERR_MUX,
    output CFG_SEND_F_ERR_MUX,
    output CFG_SYS_ERR_RC,
    output CFG_AER_RC_ERR_MUX,
    output RADM_CPL_TIMEOUT,
    output [2:0] RADM_TIMEOUT_CPL_TC,
    output [7:0] RADM_TIMEOUT_CPL_TAG,
    output [1:0] RADM_TIMEOUT_CPL_ATTR,
    output [10:0] RADM_TIMEOUT_CPL_LEN,
    output [2:0] CFG_MAX_RD_REQ_SIZE,
    output CFG_BUS_MASTER_EN,
    output [2:0] CFG_MAX_PAYLOAD_SIZE,
    output CFG_RCB,
    output CFG_MEM_SPACE_EN,
    output CFG_PM_NO_SOFT_RST,
    output CFG_CRS_SW_VIS_EN,
    output CFG_NO_SNOOP_EN,
    output CFG_RELAX_ORDER_EN,
    output [1:0] CFG_TPH_REQ_EN,
    output [2:0] CFG_PF_TPH_ST_MODE,
    output [7:0] CFG_PBUS_NUM,
    output [4:0] CFG_PBUS_DEV_NUM,
    output RBAR_CTRL_UPDATE,
    output CFG_ATOMIC_REQ_EN,
    output CFG_ATOMIC_EGRESS_BLOCK,
    output CFG_EXT_TAG_EN,
    output RADM_IDLE,
    output RADM_Q_NOT_EMPTY,
    output RADM_QOVERFLOW,
    input [1:0] DIAG_CTRL_BUS,
    input [3:0] DYN_DEBUG_INFO_SEL,
    output CFG_LINK_AUTO_BW_MUX,
    output CFG_BW_MGT_MUX,
    output CFG_PME_MUX,
    output [132:0] DEBUG_INFO_MUX,
    input APP_RAS_DES_SD_HOLD_LTSSM,
    input [1:0] APP_RAS_DES_TBA_CTRL,
    output CFG_IDO_REQ_EN,
    output CFG_IDO_CPL_EN,
    output [7:0] XADM_PH_CDTS,
    output [11:0] XADM_PD_CDTS,
    output [7:0] XADM_NPH_CDTS,
    output [11:0] XADM_NPD_CDTS,
    output [7:0] XADM_CPLH_CDTS,
    output [11:0] XADM_CPLD_CDTS,
    output [1:0] MAC_PHY_POWERDOWN,
    input [3:0] PHY_MAC_RXELECIDLE,
    input [3:0] PHY_MAC_PHYSTATUS,
    input [127:0] PHY_MAC_RXDATA,
    input [15:0] PHY_MAC_RXDATAK,
    input [3:0] PHY_MAC_RXVALID,
    input [11:0] PHY_MAC_RXSTATUS,
    output [127:0] MAC_PHY_TXDATA,
    output [15:0] MAC_PHY_TXDATAK,
    output [3:0] MAC_PHY_TXDETECTRX_LOOPBACK,
    output [3:0] MAC_PHY_TXELECIDLE_L,
    output [3:0] MAC_PHY_TXELECIDLE_H,
    output [3:0] MAC_PHY_TXCOMPLIANCE,
    output [3:0] MAC_PHY_RXPOLARITY,
    output MAC_PHY_RATE,
    output [1:0] MAC_PHY_TXDEEMPH,
    output [2:0] MAC_PHY_TXMARGIN,
    output MAC_PHY_TXSWING,
    output CFG_HW_AUTO_SP_DIS,
    input [65:0] P_DATAQ_DATAOUT,
    output [9:0] P_DATAQ_ADDRA,
    output [9:0] P_DATAQ_ADDRB,
    output [65:0] P_DATAQ_DATAIN,
    output P_DATAQ_ENA,
    output P_DATAQ_ENB,
    output P_DATAQ_WEA,
    output [10:0] XDLH_RETRYRAM_ADDR,
    output [67:0] XDLH_RETRYRAM_DATA,
    output XDLH_RETRYRAM_WE,
    output XDLH_RETRYRAM_EN,
    input [67:0] RETRYRAM_XDLH_DATA,
    output [8:0] P_HDRQ_ADDRA,
    output [8:0] P_HDRQ_ADDRB,
    output [137:0] P_HDRQ_DATAIN,
    output P_HDRQ_ENA,
    output P_HDRQ_ENB,
    output P_HDRQ_WEA,
    input [137:0] P_HDRQ_DATAOUT,
    input RAM_TEST_EN,
    input RAM_TEST_ADDRH,
    input RETRY_TEST_DATA_EN,
    input RAM_TEST_MODE_N
)  ;
endmodule


module GTP_PCIEGEN2_DFT
#(
    parameter GRS_EN = "TRUE",
    parameter PIN_MUX_INT_FORCE_EN = "FALSE",
    parameter PIN_MUX_INT_DISABLE = "FALSE",
    parameter DIAG_CTRL_BUS_B2 = "NORMAL",
    parameter DYN_DEBUG_SEL_EN = "FALSE",
    parameter integer DEBUG_INFO_SEL = 0,
    parameter integer BAR_RESIZABLE = 21,
    parameter integer NUM_OF_RBARS = 3,
    parameter integer BAR_INDEX_0 = 0,
    parameter integer BAR_INDEX_1 = 2,
    parameter integer BAR_INDEX_2 = 4,
    parameter TPH_DISABLE = "FALSE",
    parameter MSIX_CAP_DISABLE = "FALSE",
    parameter MSI_CAP_DISABLE = "FALSE",
    parameter MSI_PVM_DISABLE = "FALSE",
    parameter integer BAR_MASK_WRITABLE = 32,
    parameter integer APP_DEV_NUM = 0,
    parameter integer APP_BUS_NUM = 0,
    parameter RAM_MUX_EN = "FALSE",
    parameter ATOMIC_DISABLE = "FALSE"
) (
    input MEM_CLK,
    input PCLK,
    input PCLK_DIV2,
    input BUTTON_RST,
    input POWER_UP_RST,
    input PERST,
    output CORE_RST_N,
    output TRAINING_RST_N,
    input APP_INIT_RST,
    output PHY_RST_N,
    input [2:0] DEVICE_TYPE,
    input RX_LANE_FLIP_EN,
    input TX_LANE_FLIP_EN,
    input APP_LTSSM_EN,
    output SMLH_LINK_UP,
    output RDLH_LINK_UP,
    input APP_REQ_RETRY_EN,
    output [4:0] SMLH_LTSSM_STATE,
    output AXIS_MASTER_TVALID,
    input AXIS_MASTER_TREADY,
    output [127:0] AXIS_MASTER_TDATA,
    output [3:0] AXIS_MASTER_TKEEP,
    output AXIS_MASTER_TLAST,
    output [7:0] AXIS_MASTER_TUSER,
    input [2:0] TRGT1_RADM_PKT_HALT,
    output [5:0] RADM_GRANT_TLP_TYPE,
    output AXIS_SLAVE0_TREADY,
    input AXIS_SLAVE0_TVALID,
    input [127:0] AXIS_SLAVE0_TDATA,
    input AXIS_SLAVE0_TLAST,
    input AXIS_SLAVE0_TUSER,
    output AXIS_SLAVE1_TREADY,
    input AXIS_SLAVE1_TVALID,
    input [127:0] AXIS_SLAVE1_TDATA,
    input AXIS_SLAVE1_TLAST,
    input AXIS_SLAVE1_TUSER,
    output AXIS_SLAVE2_TREADY,
    input AXIS_SLAVE2_TVALID,
    input [127:0] AXIS_SLAVE2_TDATA,
    input AXIS_SLAVE2_TLAST,
    input AXIS_SLAVE2_TUSER,
    output PM_XTLH_BLOCK_TLP,
    input [31:0] DBI_ADDR,
    input [31:0] DBI_DIN,
    input DBI_CS,
    input DBI_CS2,
    input [3:0] DBI_WR,
    input APP_DBI_RO_WR_DISABLE,
    output LBC_DBI_ACK,
    output [31:0] LBC_DBI_DOUT,
    output SEDO,
    output SEDO_EN,
    input SEDI,
    input SEDI_ACK,
    output CFG_INT_DISABLE,
    input SYS_INT,
    output INTA_GRT_MUX,
    output INTB_GRT_MUX,
    output INTC_GRT_MUX,
    output INTD_GRT_MUX,
    input VEN_MSI_REQ,
    input [2:0] VEN_MSI_TC,
    input [4:0] VEN_MSI_VECTOR,
    output VEN_MSI_GRANT,
    input [31:0] CFG_MSI_PENDING,
    output CFG_MSI_EN,
    input [63:0] MSIX_ADDR,
    input [31:0] MSIX_DATA,
    output CFG_MSIX_EN,
    output CFG_MSIX_FUNC_MASK,
    output RADM_PM_TURNOFF,
    output RADM_MSG_UNLOCK,
    input OUTBAND_PWRUP_CMD,
    output PM_STATUS,
    output [2:0] PM_DSTATE,
    output AUX_PM_EN,
    output PM_PME_EN,
    output PM_LINKST_IN_L0S,
    output PM_LINKST_IN_L1,
    output PM_LINKST_IN_L2,
    output PM_LINKST_L2_EXIT,
    input APP_REQ_ENTR_L1,
    input APP_READY_ENTR_L23,
    input APP_REQ_EXIT_L1,
    input APP_XFER_PENDING,
    output WAKE,
    output RADM_PM_PME,
    output RADM_PM_TO_ACK,
    input APPS_PM_XMT_TURNOFF,
    input APP_UNLOCK_MSG,
    input APPS_PM_XMT_PME,
    input APP_CLK_PM_EN,
    output [4:0] PM_MASTER_STATE,
    output [4:0] PM_SLAVE_STATE,
    input SYS_AUX_PWR_DET,
    input APP_HDR_VALID,
    input [127:0] APP_HDR_LOG,
    input [12:0] APP_ERR_BUS,
    input APP_ERR_ADVISORY,
    output CFG_SEND_COR_ERR_MUX,
    output CFG_SEND_NF_ERR_MUX,
    output CFG_SEND_F_ERR_MUX,
    output CFG_SYS_ERR_RC,
    output CFG_AER_RC_ERR_MUX,
    output RADM_CPL_TIMEOUT,
    output [2:0] RADM_TIMEOUT_CPL_TC,
    output [7:0] RADM_TIMEOUT_CPL_TAG,
    output [1:0] RADM_TIMEOUT_CPL_ATTR,
    output [10:0] RADM_TIMEOUT_CPL_LEN,
    output [2:0] CFG_MAX_RD_REQ_SIZE,
    output CFG_BUS_MASTER_EN,
    output [2:0] CFG_MAX_PAYLOAD_SIZE,
    output CFG_RCB,
    output CFG_MEM_SPACE_EN,
    output CFG_PM_NO_SOFT_RST,
    output CFG_CRS_SW_VIS_EN,
    output CFG_NO_SNOOP_EN,
    output CFG_RELAX_ORDER_EN,
    output [1:0] CFG_TPH_REQ_EN,
    output [2:0] CFG_PF_TPH_ST_MODE,
    output [7:0] CFG_PBUS_NUM,
    output [4:0] CFG_PBUS_DEV_NUM,
    output RBAR_CTRL_UPDATE,
    output CFG_ATOMIC_REQ_EN,
    output CFG_ATOMIC_EGRESS_BLOCK,
    output CFG_EXT_TAG_EN,
    output RADM_IDLE,
    output RADM_Q_NOT_EMPTY,
    output RADM_QOVERFLOW,
    input [1:0] DIAG_CTRL_BUS,
    input [3:0] DYN_DEBUG_INFO_SEL,
    output CFG_LINK_AUTO_BW_MUX,
    output CFG_BW_MGT_MUX,
    output CFG_PME_MUX,
    output [132:0] DEBUG_INFO_MUX,
    input APP_RAS_DES_SD_HOLD_LTSSM,
    input [1:0] APP_RAS_DES_TBA_CTRL,
    output CFG_IDO_REQ_EN,
    output CFG_IDO_CPL_EN,
    output [7:0] XADM_PH_CDTS,
    output [11:0] XADM_PD_CDTS,
    output [7:0] XADM_NPH_CDTS,
    output [11:0] XADM_NPD_CDTS,
    output [7:0] XADM_CPLH_CDTS,
    output [11:0] XADM_CPLD_CDTS,
    output [1:0] MAC_PHY_POWERDOWN,
    input [3:0] PHY_MAC_RXELECIDLE,
    input [3:0] PHY_MAC_PHYSTATUS,
    input [127:0] PHY_MAC_RXDATA,
    input [15:0] PHY_MAC_RXDATAK,
    input [3:0] PHY_MAC_RXVALID,
    input [11:0] PHY_MAC_RXSTATUS,
    output [127:0] MAC_PHY_TXDATA,
    output [15:0] MAC_PHY_TXDATAK,
    output [3:0] MAC_PHY_TXDETECTRX_LOOPBACK,
    output [3:0] MAC_PHY_TXELECIDLE_L,
    output [3:0] MAC_PHY_TXELECIDLE_H,
    output [3:0] MAC_PHY_TXCOMPLIANCE,
    output [3:0] MAC_PHY_RXPOLARITY,
    output MAC_PHY_RATE,
    output [1:0] MAC_PHY_TXDEEMPH,
    output [2:0] MAC_PHY_TXMARGIN,
    output MAC_PHY_TXSWING,
    output CFG_HW_AUTO_SP_DIS,
    input [65:0] P_DATAQ_DATAOUT,
    output [9:0] P_DATAQ_ADDRA,
    output [9:0] P_DATAQ_ADDRB,
    output [65:0] P_DATAQ_DATAIN,
    output P_DATAQ_ENA,
    output P_DATAQ_ENB,
    output P_DATAQ_WEA,
    output [10:0] XDLH_RETRYRAM_ADDR,
    output [67:0] XDLH_RETRYRAM_DATA,
    output XDLH_RETRYRAM_WE,
    output XDLH_RETRYRAM_EN,
    input [67:0] RETRYRAM_XDLH_DATA,
    output [8:0] P_HDRQ_ADDRA,
    output [8:0] P_HDRQ_ADDRB,
    output [137:0] P_HDRQ_DATAIN,
    output P_HDRQ_ENA,
    output P_HDRQ_ENB,
    output P_HDRQ_WEA,
    input [137:0] P_HDRQ_DATAOUT,
    input RAM_TEST_EN,
    input RAM_TEST_ADDRH,
    input RETRY_TEST_DATA_EN,
    input RAM_TEST_MODE_N,
    input TEST_SE_N,
    input TEST_RST_N,
    input TEST_MODE_N
)  ;
endmodule


module GTP_PCIEGEN3
#(
    parameter PF1_ENABLE = "TRUE",
    parameter FLT_SHORT_TLP = "TRUE",
    parameter integer APP_DEV_NUM = 0,
    parameter integer APP_BUS_NUM = 0,
    parameter integer DEBUG_INFO_SEL = 0,
    parameter DYN_DEBUG_SEL_EN = "FALSE",
    parameter GRS_EN = "FALSE",
    parameter VF_ER_REPORT_EN = "TRUE",
    parameter ATOMIC_DISABLE = "FALSE",
    parameter VC_DISABLE = "FALSE",
    parameter SRIOV_DISABLE = "FALSE",
    parameter integer BAR_RESIZABLE = 1365,
    parameter integer NUM_OF_RBARS = 27,
    parameter integer MSI_PVM_DISABLE = 0,
    parameter integer BAR_MASK_WRITABLE = 0
) (
    input PCLK,
    input PCLK_DIV2,
    input MEM_CLK,
    input USER_CLK,
    input BUTTON_RST,
    input POWER_UP_RST,
    input PERST,
    output USER_RST_N,
    output TRAINING_RST_N,
    input APP_INIT_RST,
    output PHY_RST_N,
    input [3:0] DEVICE_TYPE,
    input RX_LANE_FLIP_EN,
    input TX_LANE_FLIP_EN,
    input APP_LTSSM_ENABLE,
    output SMLH_LINK_UP,
    output RDLH_LINK_UP,
    input APP_REQ_RETRY_EN,
    output [5:0] SMLH_LTSSM_STATE,
    output CFG_2ND_RESET,
    output LINK_REQ_RST,
    input [1:0] APP_PF_REQ_RETRY_EN,
    output [5:0] CFG_VF_BME,
    input [5:0] APP_VF_REQ_RETRY_EN,
    output SMLH_REQ_RST,
    output [255:0] AXIS_MASTER0_TDATA,
    output [7:0] AXIS_MASTER0_TKEEP,
    output AXIS_MASTER0_TLAST,
    output [12:0] AXIS_MASTER0_TUSER,
    output AXIS_MASTER0_TVALID,
    input AXIS_MASTER0_TREADY,
    input USER_RCVD_NP_READY,
    output [5:0] CORE_AVL_NP_CNT,
    input USER_RCVD_P_READY,
    output [5:0] CORE_AVL_P_CNT,
    output [255:0] AXIS_MASTER1_TDATA,
    output [7:0] AXIS_MASTER1_TKEEP,
    output [33:0] AXIS_MASTER1_TUSER,
    output AXIS_MASTER1_TVALID,
    input [255:0] AXIS_SLAVE0_TDATA,
    input AXIS_SLAVE0_TLAST,
    input [5:0] AXIS_SLAVE0_TUSER,
    input AXIS_SLAVE0_TVALID,
    output AXIS_SLAVE0_TREADY,
    input [255:0] AXIS_SLAVE1_TDATA,
    input AXIS_SLAVE1_TLAST,
    input [5:0] AXIS_SLAVE1_TUSER,
    input AXIS_SLAVE1_TVALID,
    output AXIS_SLAVE1_TREADY,
    input [255:0] AXIS_SLAVE2_TDATA,
    input AXIS_SLAVE2_TLAST,
    input [5:0] AXIS_SLAVE2_TUSER,
    input AXIS_SLAVE2_TVALID,
    output AXIS_SLAVE2_TREADY,
    output [1:0] RADM_CPL_TIMEOUT,
    output [3:0] RADM_TIMEOUT_CPL_ATTR,
    output [21:0] RADM_TIMEOUT_CPL_LEN,
    output [15:0] RADM_TIMEOUT_CPL_TAG,
    output [5:0] RADM_TIMEOUT_CPL_TC,
    output [1:0] RADM_TIMEOUT_FUNC_NUM,
    output [1:0] RADM_TIMEOUT_VFUNC_ACTIVE,
    output [5:0] RADM_TIMEOUT_VFUNC_NUM,
    input APP_DBI_RO_WR_DISABLE,
    input [31:0] DBI_ADDR,
    input DBI_CS,
    input DBI_CS2,
    input [31:0] DBI_DIN,
    input DBI_FUNC_NUM,
    input DBI_VFUNC_ACTIVE,
    input [2:0] DBI_VFUNC_NUM,
    input [3:0] DBI_WR,
    output LBC_DBI_ACK,
    output [31:0] LBC_DBI_DOUT,
    input [1:0] SEDI,
    input [1:0] SEDI_ACK,
    output [1:0] SEDO,
    output [1:0] SEDO_EN,
    input [1:0] SYS_INT,
    output [1:0] CFG_INT_DISABLE,
    output INT_GRT,
    input [63:0] CFG_MSI_PENDING,
    input [191:0] CFG_VF_MSI_PENDING,
    input VEN_MSI_FUNC_NUM,
    input VEN_MSI_REQ,
    input [2:0] VEN_MSI_TC,
    input [4:0] VEN_MSI_VECTOR,
    input VEN_MSI_VFUNC_ACTIVE,
    input [2:0] VEN_MSI_VFUNC_NUM,
    output [1:0] CFG_MSI_EN,
    output CFG_MSI_MASK_UPDATE,
    output [5:0] CFG_MULTI_MSI_EN,
    output [5:0] CFG_VF_MSI_EN,
    output [17:0] CFG_VF_MULTI_MSI_EN,
    output VEN_MSI_GRANT,
    input [63:0] MSIX_ADDR,
    input [31:0] MSIX_DATA,
    output [1:0] CFG_MSIX_EN,
    output [1:0] CFG_MSIX_FUNC_MASK,
    output [5:0] CFG_VF_MSIX_EN,
    output [5:0] CFG_VF_MSIX_FUNC_MASK,
    output CFG_BW_MGT_MSI,
    output CFG_LINK_AUTO_BW_MSI,
    output [1:0] CFG_PME_MSI,
    output CFG_BW_MGT_INT,
    output CFG_LINK_AUTO_BW_INT,
    output CFG_LINK_EQ_REQ_INT,
    output [1:0] CFG_PME_INT,
    output [1:0] CFG_NF_ERR_RPT_EN,
    output [1:0] CFG_NO_SNOOP_EN,
    output [1:0] CFG_OBFF_EN,
    output [4:0] CFG_PBUS_DEV_NUM,
    output [7:0] CFG_PBUS_NUM,
    output [1:0] CFG_MEM_SPACE_EN,
    output [1:0] CFG_EXT_TAG_EN,
    output [1:0] CFG_F_ERR_RPT_EN,
    output [1:0] CFG_ARI_FWD_EN,
    output [1:0] CFG_ATOMIC_EGRESS_BLOCK,
    output [1:0] CFG_ATOMIC_REQ_EN,
    output [1:0] CFG_BUS_MASTER_EN,
    output [1:0] CFG_COR_ERR_RPT_EN,
    output [1:0] CFG_CRS_SW_VIS_EN,
    output [5:0] CFG_MAX_PAYLOAD_SIZE,
    output [5:0] CFG_MAX_RD_REQ_SIZE,
    output [1:0] CFG_VF_EN,
    output [7:0] CFG_TC_ENABLE,
    output [1:0] CFG_RCB,
    output [1:0] CFG_REG_SERREN,
    output [1:0] CFG_RELAX_ORDER_EN,
    output [1:0] RBAR_CTRL_UPDATE,
    input APP_CLK_PM_EN,
    input [5:0] APPS_PM_VF_XMT_PME,
    input [1:0] APPS_PM_XMT_PME,
    input APPS_PM_XMT_TURNOFF,
    input APP_UNLOCK_MSG,
    output [1:0] AUX_PM_EN,
    output [5:0] PM_DSTATE,
    output [4:0] PM_MASTER_STATE,
    output [1:0] PM_PME_EN,
    output [4:0] PM_SLAVE_STATE,
    output [1:0] PM_STATUS,
    output [17:0] PM_VF_DSTATE,
    output [5:0] PM_VF_PME_EN,
    output [5:0] PM_VF_STATUS,
    output PM_XTLH_BLOCK_TLP,
    input APP_READY_ENTR_L23,
    input APP_REQ_ENTR_L1,
    input APP_REQ_EXIT_L1,
    input [31:0] CFG_PWR_BUDGET_DATA_REG,
    input CFG_PWR_BUDGET_FUNC_NUM,
    input CFG_PWR_BUDGET_VALID,
    output [1:0] DPA_SUBSTATE_UPDATE,
    output WAKE,
    output [7:0] CFG_PWR_BUDGET_DATA_SEL_REG,
    output [1:0] CFG_PWR_BUDGET_SEL,
    input APP_XFER_PENDING,
    input [127:0] APP_HDR_LOG,
    input APP_HDR_VALID,
    input APP_ERR_ADVISORY,
    input [12:0] APP_ERR_BUS,
    input APP_ERR_FUNC_NUM,
    input APP_ERR_VFUNC_ACTIVE,
    input [2:0] APP_ERR_VFUNC_NUM,
    output [1:0] CFG_SEND_COR_ERR,
    output [1:0] CFG_SEND_F_ERR,
    output [1:0] CFG_SEND_NF_ERR,
    output [1:0] CFG_AER_RC_ERR_INT,
    output [1:0] CFG_AER_RC_ERR_MSI,
    output [1:0] CFG_SYS_ERR_RC,
    input APP_LTR_MSG_FUNC_NUM,
    input [31:0] APP_LTR_MSG_LATENCY,
    input APP_LTR_MSG_REQ,
    output APP_LTR_MSG_GRANT,
    output CFG_LTR_M_EN,
    output CFG_DISABLE_LTR_CLR_MSG,
    input [1:0] APP_FLR_PF_DONE,
    input [5:0] APP_FLR_VF_DONE,
    output [1:0] CFG_FLR_PF_ACTIVE,
    output [5:0] CFG_FLR_VF_ACTIVE,
    output [5:0] CFG_START_VFI,
    output [5:0] CFG_NUM_VF,
    input APP_OBFF_CPU_ACTIVE_MSG_REQ,
    input APP_OBFF_IDLE_MSG_REQ,
    input APP_OBFF_OBFF_MSG_REQ,
    output APP_OBFF_MSG_GRANT,
    output MSG_RCVD,
    output [7:0] MSG_RCVD_DATA,
    output [4:0] MSG_RCVD_TYPE,
    input APP_RAS_DES_SD_HOLD_LTSSM,
    input [2:0] DIAG_CTRL_BUS,
    input [5:0] DYN_DEBUG_INFO_SEL,
    output [142:0] DEBUG_INFO_MUX,
    output [1:0] CFG_IDO_CPL_EN,
    output [1:0] CFG_IDO_REQ_EN,
    output [11:0] XADM_CPLD_CDTS,
    output [7:0] XADM_CPLH_CDTS,
    output [11:0] XADM_NPD_CDTS,
    output [7:0] XADM_NPH_CDTS,
    output [11:0] XADM_PD_CDTS,
    output [7:0] XADM_PH_CDTS,
    output RADM_Q_NOT_EMPTY,
    output RADM_QOVERFLOW,
    input [47:0] PHY_MAC_DIRFEEDBACK,
    input [63:0] PHY_MAC_FOMFEEDBACK,
    input [47:0] PHY_MAC_LOCALFS,
    input [47:0] PHY_MAC_LOCALLF,
    input [7:0] PHY_MAC_LOCAL_TX_COEF_VALID,
    input [47:0] PHY_MAC_LOCAL_TX_PSET_COEF,
    input [7:0] PHY_MAC_PHYSTATUS,
    input [255:0] PHY_MAC_RXDATA,
    input [31:0] PHY_MAC_RXDATAK,
    input [7:0] PHY_MAC_RXDATAVALID,
    input [7:0] PHY_MAC_RXELECIDLE,
    input [7:0] PHY_MAC_RXSTARTBLOCK,
    input [23:0] PHY_MAC_RXSTATUS,
    input [15:0] PHY_MAC_RXSYNCHEADER,
    input [7:0] PHY_MAC_RXVALID,
    output MAC_PHY_BLOCKALIGNCONTROL,
    output [7:0] MAC_PHY_DIRCHANGE,
    output [47:0] MAC_PHY_FS,
    output [7:0] MAC_PHY_GETLOCAL_PSET_COEF,
    output [7:0] MAC_PHY_INVALID_REQ,
    output [47:0] MAC_PHY_LF,
    output [31:0] MAC_PHY_LOCAL_PSET_INDEX,
    output [1:0] MAC_PHY_POWERDOWN,
    output [1:0] MAC_PHY_RATE,
    output [7:0] MAC_PHY_RXEQEVAL,
    output [7:0] MAC_PHY_RXEQINPROGRESS,
    output [7:0] MAC_PHY_RXPOLARITY,
    output [23:0] MAC_PHY_RXPRESETHINT,
    output [7:0] MAC_PHY_TXCOMPLIANCE,
    output [255:0] MAC_PHY_TXDATA,
    output [31:0] MAC_PHY_TXDATAK,
    output [7:0] MAC_PHY_TXDATAVALID,
    output [48:0] MAC_PHY_TXDEEMPH,
    output [7:0] MAC_PHY_TXDETECTRX_LOOPBACK,
    output [7:0] MAC_PHY_TXELECIDLE_H,
    output [7:0] MAC_PHY_TXELECIDLE_L,
    output [2:0] MAC_PHY_TXMARGIN,
    output [7:0] MAC_PHY_TXSTARTBLOCK,
    output MAC_PHY_TXSWING,
    output [15:0] MAC_PHY_TXSYNCHEADER,
    output [9:0] PNP_RAM_RD_ADDR,
    output PNP_RAM_RD_EN,
    output [9:0] PNP_RAM_WR_ADDR,
    output [134:0] PNP_RAM_WR_DATA,
    output PNP_RAM_WR_EN,
    input [134:0] PNP_RAM_RD_DATA,
    input [134:0] RETRYRAM_XDLH_DATA,
    output [9:0] XDLH_RETRYRAM_ADDR,
    output [134:0] XDLH_RETRYRAM_DATA,
    output XDLH_RETRYRAM_EN,
    output XDLH_RETRYRAM_WE,
    output [5:0] CFG_PF_TPH_ST_MODE,
    output [1:0] CFG_TPH_REQ_EN,
    output [5:0] CFG_VF_TPH_REQ_EN,
    output [17:0] CFG_VF_TPH_ST_MODE,
    input TPH_RD_DATA_VALID,
    input [15:0] TPH_RAM_RD_DATA,
    output [4:0] TPH_RAM_ADDR,
    output [2:0] TPH_RAM_FUNC_NUM,
    output TPH_RAM_FUNC_ACTIVE,
    output [1:0] TPH_RAM_WR_BYTE_EN,
    output [15:0] TPH_RAM_WR_DATA,
    output TPH_RAM_WR_EN,
    input RAM_TEST_EN,
    input RAM_TEST_ADDRH,
    input RETRY_TEST_DATA_EN,
    input RAM_TEST_MODE_N
)  ;
endmodule


module GTP_PCIEGEN3_DFT
#(
    parameter PF1_ENABLE = "TRUE",
    parameter FLT_SHORT_TLP = "TRUE",
    parameter integer APP_DEV_NUM = 0,
    parameter integer APP_BUS_NUM = 0,
    parameter integer DEBUG_INFO_SEL = 0,
    parameter DYN_DEBUG_SEL_EN = "FALSE",
    parameter GRS_EN = "FALSE",
    parameter VF_ER_REPORT_EN = "TRUE",
    parameter ATOMIC_DISABLE = "FALSE",
    parameter VC_DISABLE = "FALSE",
    parameter SRIOV_DISABLE = "FALSE",
    parameter integer BAR_RESIZABLE = 1365,
    parameter integer NUM_OF_RBARS = 27,
    parameter integer MSI_PVM_DISABLE = 0,
    parameter integer BAR_MASK_WRITABLE = 0
) (
    input PCLK,
    input PCLK_DIV2,
    input MEM_CLK,
    input USER_CLK,
    input BUTTON_RST,
    input POWER_UP_RST,
    input PERST,
    output USER_RST_N,
    output TRAINING_RST_N,
    input APP_INIT_RST,
    output PHY_RST_N,
    input [3:0] DEVICE_TYPE,
    input RX_LANE_FLIP_EN,
    input TX_LANE_FLIP_EN,
    input APP_LTSSM_ENABLE,
    output SMLH_LINK_UP,
    output RDLH_LINK_UP,
    input APP_REQ_RETRY_EN,
    output [5:0] SMLH_LTSSM_STATE,
    output CFG_2ND_RESET,
    output LINK_REQ_RST,
    input [1:0] APP_PF_REQ_RETRY_EN,
    output [5:0] CFG_VF_BME,
    input [5:0] APP_VF_REQ_RETRY_EN,
    output SMLH_REQ_RST,
    output [255:0] AXIS_MASTER0_TDATA,
    output [7:0] AXIS_MASTER0_TKEEP,
    output AXIS_MASTER0_TLAST,
    output [12:0] AXIS_MASTER0_TUSER,
    output AXIS_MASTER0_TVALID,
    input AXIS_MASTER0_TREADY,
    input USER_RCVD_NP_READY,
    output [5:0] CORE_AVL_NP_CNT,
    input USER_RCVD_P_READY,
    output [5:0] CORE_AVL_P_CNT,
    output [255:0] AXIS_MASTER1_TDATA,
    output [7:0] AXIS_MASTER1_TKEEP,
    output [33:0] AXIS_MASTER1_TUSER,
    output AXIS_MASTER1_TVALID,
    input [255:0] AXIS_SLAVE0_TDATA,
    input AXIS_SLAVE0_TLAST,
    input [5:0] AXIS_SLAVE0_TUSER,
    input AXIS_SLAVE0_TVALID,
    output AXIS_SLAVE0_TREADY,
    input [255:0] AXIS_SLAVE1_TDATA,
    input AXIS_SLAVE1_TLAST,
    input [5:0] AXIS_SLAVE1_TUSER,
    input AXIS_SLAVE1_TVALID,
    output AXIS_SLAVE1_TREADY,
    input [255:0] AXIS_SLAVE2_TDATA,
    input AXIS_SLAVE2_TLAST,
    input [5:0] AXIS_SLAVE2_TUSER,
    input AXIS_SLAVE2_TVALID,
    output AXIS_SLAVE2_TREADY,
    output [1:0] RADM_CPL_TIMEOUT,
    output [3:0] RADM_TIMEOUT_CPL_ATTR,
    output [21:0] RADM_TIMEOUT_CPL_LEN,
    output [15:0] RADM_TIMEOUT_CPL_TAG,
    output [5:0] RADM_TIMEOUT_CPL_TC,
    output [1:0] RADM_TIMEOUT_FUNC_NUM,
    output [1:0] RADM_TIMEOUT_VFUNC_ACTIVE,
    output [5:0] RADM_TIMEOUT_VFUNC_NUM,
    input APP_DBI_RO_WR_DISABLE,
    input [31:0] DBI_ADDR,
    input DBI_CS,
    input DBI_CS2,
    input [31:0] DBI_DIN,
    input DBI_FUNC_NUM,
    input DBI_VFUNC_ACTIVE,
    input [2:0] DBI_VFUNC_NUM,
    input [3:0] DBI_WR,
    output LBC_DBI_ACK,
    output [31:0] LBC_DBI_DOUT,
    input [1:0] SEDI,
    input [1:0] SEDI_ACK,
    output [1:0] SEDO,
    output [1:0] SEDO_EN,
    input [1:0] SYS_INT,
    output [1:0] CFG_INT_DISABLE,
    output INT_GRT,
    input [63:0] CFG_MSI_PENDING,
    input [191:0] CFG_VF_MSI_PENDING,
    input VEN_MSI_FUNC_NUM,
    input VEN_MSI_REQ,
    input [2:0] VEN_MSI_TC,
    input [4:0] VEN_MSI_VECTOR,
    input VEN_MSI_VFUNC_ACTIVE,
    input [2:0] VEN_MSI_VFUNC_NUM,
    output [1:0] CFG_MSI_EN,
    output CFG_MSI_MASK_UPDATE,
    output [5:0] CFG_MULTI_MSI_EN,
    output [5:0] CFG_VF_MSI_EN,
    output [17:0] CFG_VF_MULTI_MSI_EN,
    output VEN_MSI_GRANT,
    input [63:0] MSIX_ADDR,
    input [31:0] MSIX_DATA,
    output [1:0] CFG_MSIX_EN,
    output [1:0] CFG_MSIX_FUNC_MASK,
    output [5:0] CFG_VF_MSIX_EN,
    output [5:0] CFG_VF_MSIX_FUNC_MASK,
    output CFG_BW_MGT_MSI,
    output CFG_LINK_AUTO_BW_MSI,
    output [1:0] CFG_PME_MSI,
    output CFG_BW_MGT_INT,
    output CFG_LINK_AUTO_BW_INT,
    output CFG_LINK_EQ_REQ_INT,
    output [1:0] CFG_PME_INT,
    output [1:0] CFG_NF_ERR_RPT_EN,
    output [1:0] CFG_NO_SNOOP_EN,
    output [1:0] CFG_OBFF_EN,
    output [4:0] CFG_PBUS_DEV_NUM,
    output [7:0] CFG_PBUS_NUM,
    output [1:0] CFG_MEM_SPACE_EN,
    output [1:0] CFG_EXT_TAG_EN,
    output [1:0] CFG_F_ERR_RPT_EN,
    output [1:0] CFG_ARI_FWD_EN,
    output [1:0] CFG_ATOMIC_EGRESS_BLOCK,
    output [1:0] CFG_ATOMIC_REQ_EN,
    output [1:0] CFG_BUS_MASTER_EN,
    output [1:0] CFG_COR_ERR_RPT_EN,
    output [1:0] CFG_CRS_SW_VIS_EN,
    output [5:0] CFG_MAX_PAYLOAD_SIZE,
    output [5:0] CFG_MAX_RD_REQ_SIZE,
    output [1:0] CFG_VF_EN,
    output [7:0] CFG_TC_ENABLE,
    output [1:0] CFG_RCB,
    output [1:0] CFG_REG_SERREN,
    output [1:0] CFG_RELAX_ORDER_EN,
    output [1:0] RBAR_CTRL_UPDATE,
    input APP_CLK_PM_EN,
    input [5:0] APPS_PM_VF_XMT_PME,
    input [1:0] APPS_PM_XMT_PME,
    input APPS_PM_XMT_TURNOFF,
    input APP_UNLOCK_MSG,
    output [1:0] AUX_PM_EN,
    output [5:0] PM_DSTATE,
    output [4:0] PM_MASTER_STATE,
    output [1:0] PM_PME_EN,
    output [4:0] PM_SLAVE_STATE,
    output [1:0] PM_STATUS,
    output [17:0] PM_VF_DSTATE,
    output [5:0] PM_VF_PME_EN,
    output [5:0] PM_VF_STATUS,
    output PM_XTLH_BLOCK_TLP,
    input APP_READY_ENTR_L23,
    input APP_REQ_ENTR_L1,
    input APP_REQ_EXIT_L1,
    input [31:0] CFG_PWR_BUDGET_DATA_REG,
    input CFG_PWR_BUDGET_FUNC_NUM,
    input CFG_PWR_BUDGET_VALID,
    output [1:0] DPA_SUBSTATE_UPDATE,
    output WAKE,
    output [7:0] CFG_PWR_BUDGET_DATA_SEL_REG,
    output [1:0] CFG_PWR_BUDGET_SEL,
    input APP_XFER_PENDING,
    input [127:0] APP_HDR_LOG,
    input APP_HDR_VALID,
    input APP_ERR_ADVISORY,
    input [12:0] APP_ERR_BUS,
    input APP_ERR_FUNC_NUM,
    input APP_ERR_VFUNC_ACTIVE,
    input [2:0] APP_ERR_VFUNC_NUM,
    output [1:0] CFG_SEND_COR_ERR,
    output [1:0] CFG_SEND_F_ERR,
    output [1:0] CFG_SEND_NF_ERR,
    output [1:0] CFG_AER_RC_ERR_INT,
    output [1:0] CFG_AER_RC_ERR_MSI,
    output [1:0] CFG_SYS_ERR_RC,
    input APP_LTR_MSG_FUNC_NUM,
    input [31:0] APP_LTR_MSG_LATENCY,
    input APP_LTR_MSG_REQ,
    output APP_LTR_MSG_GRANT,
    output CFG_LTR_M_EN,
    output CFG_DISABLE_LTR_CLR_MSG,
    input [1:0] APP_FLR_PF_DONE,
    input [5:0] APP_FLR_VF_DONE,
    output [1:0] CFG_FLR_PF_ACTIVE,
    output [5:0] CFG_FLR_VF_ACTIVE,
    output [5:0] CFG_START_VFI,
    output [5:0] CFG_NUM_VF,
    input APP_OBFF_CPU_ACTIVE_MSG_REQ,
    input APP_OBFF_IDLE_MSG_REQ,
    input APP_OBFF_OBFF_MSG_REQ,
    output APP_OBFF_MSG_GRANT,
    output MSG_RCVD,
    output [7:0] MSG_RCVD_DATA,
    output [4:0] MSG_RCVD_TYPE,
    input APP_RAS_DES_SD_HOLD_LTSSM,
    input [2:0] DIAG_CTRL_BUS,
    input [5:0] DYN_DEBUG_INFO_SEL,
    output [142:0] DEBUG_INFO_MUX,
    output [1:0] CFG_IDO_CPL_EN,
    output [1:0] CFG_IDO_REQ_EN,
    output [11:0] XADM_CPLD_CDTS,
    output [7:0] XADM_CPLH_CDTS,
    output [11:0] XADM_NPD_CDTS,
    output [7:0] XADM_NPH_CDTS,
    output [11:0] XADM_PD_CDTS,
    output [7:0] XADM_PH_CDTS,
    output RADM_Q_NOT_EMPTY,
    output RADM_QOVERFLOW,
    input [47:0] PHY_MAC_DIRFEEDBACK,
    input [63:0] PHY_MAC_FOMFEEDBACK,
    input [47:0] PHY_MAC_LOCALFS,
    input [47:0] PHY_MAC_LOCALLF,
    input [7:0] PHY_MAC_LOCAL_TX_COEF_VALID,
    input [47:0] PHY_MAC_LOCAL_TX_PSET_COEF,
    input [7:0] PHY_MAC_PHYSTATUS,
    input [255:0] PHY_MAC_RXDATA,
    input [31:0] PHY_MAC_RXDATAK,
    input [7:0] PHY_MAC_RXDATAVALID,
    input [7:0] PHY_MAC_RXELECIDLE,
    input [7:0] PHY_MAC_RXSTARTBLOCK,
    input [23:0] PHY_MAC_RXSTATUS,
    input [15:0] PHY_MAC_RXSYNCHEADER,
    input [7:0] PHY_MAC_RXVALID,
    output MAC_PHY_BLOCKALIGNCONTROL,
    output [7:0] MAC_PHY_DIRCHANGE,
    output [47:0] MAC_PHY_FS,
    output [7:0] MAC_PHY_GETLOCAL_PSET_COEF,
    output [7:0] MAC_PHY_INVALID_REQ,
    output [47:0] MAC_PHY_LF,
    output [31:0] MAC_PHY_LOCAL_PSET_INDEX,
    output [1:0] MAC_PHY_POWERDOWN,
    output [1:0] MAC_PHY_RATE,
    output [7:0] MAC_PHY_RXEQEVAL,
    output [7:0] MAC_PHY_RXEQINPROGRESS,
    output [7:0] MAC_PHY_RXPOLARITY,
    output [23:0] MAC_PHY_RXPRESETHINT,
    output [7:0] MAC_PHY_TXCOMPLIANCE,
    output [255:0] MAC_PHY_TXDATA,
    output [31:0] MAC_PHY_TXDATAK,
    output [7:0] MAC_PHY_TXDATAVALID,
    output [48:0] MAC_PHY_TXDEEMPH,
    output [7:0] MAC_PHY_TXDETECTRX_LOOPBACK,
    output [7:0] MAC_PHY_TXELECIDLE_H,
    output [7:0] MAC_PHY_TXELECIDLE_L,
    output [2:0] MAC_PHY_TXMARGIN,
    output [7:0] MAC_PHY_TXSTARTBLOCK,
    output MAC_PHY_TXSWING,
    output [15:0] MAC_PHY_TXSYNCHEADER,
    output [9:0] PNP_RAM_RD_ADDR,
    output PNP_RAM_RD_EN,
    output [9:0] PNP_RAM_WR_ADDR,
    output [134:0] PNP_RAM_WR_DATA,
    output PNP_RAM_WR_EN,
    input [134:0] PNP_RAM_RD_DATA,
    input [134:0] RETRYRAM_XDLH_DATA,
    output [9:0] XDLH_RETRYRAM_ADDR,
    output [134:0] XDLH_RETRYRAM_DATA,
    output XDLH_RETRYRAM_EN,
    output XDLH_RETRYRAM_WE,
    output [5:0] CFG_PF_TPH_ST_MODE,
    output [1:0] CFG_TPH_REQ_EN,
    output [5:0] CFG_VF_TPH_REQ_EN,
    output [17:0] CFG_VF_TPH_ST_MODE,
    input TPH_RD_DATA_VALID,
    input [15:0] TPH_RAM_RD_DATA,
    output [4:0] TPH_RAM_ADDR,
    output [2:0] TPH_RAM_FUNC_NUM,
    output TPH_RAM_FUNC_ACTIVE,
    output [1:0] TPH_RAM_WR_BYTE_EN,
    output [15:0] TPH_RAM_WR_DATA,
    output TPH_RAM_WR_EN,
    input RAM_TEST_EN,
    input RAM_TEST_ADDRH,
    input RETRY_TEST_DATA_EN,
    input RAM_TEST_MODE_N,
    input TEST_MODE_N,
    input TEST_RST_N,
    input TEST_SE_N
)  ;
endmodule


module GTP_PPLL
#(
    parameter real CLKIN_FREQ = 50.0,
    parameter LOCK_MODE = 1'b0,
    parameter integer STATIC_RATIOI = 1,
    parameter integer STATIC_RATIOM = 1,
    parameter integer STATIC_RATIO0 = 1,
    parameter integer STATIC_RATIO1 = 1,
    parameter integer STATIC_RATIO2 = 1,
    parameter integer STATIC_RATIO3 = 1,
    parameter integer STATIC_RATIO4 = 1,
    parameter integer STATIC_RATIOPHY = 1,
    parameter integer STATIC_RATIOF = 1,
    parameter integer STATIC_DUTY0 = 2,
    parameter integer STATIC_DUTY1 = 2,
    parameter integer STATIC_DUTY2 = 2,
    parameter integer STATIC_DUTY3 = 2,
    parameter integer STATIC_DUTY4 = 2,
    parameter integer STATIC_DUTYPHY = 2,
    parameter integer STATIC_DUTYF = 2,
    parameter integer STATIC_PHASE0 = 0,
    parameter integer STATIC_PHASE1 = 0,
    parameter integer STATIC_PHASE2 = 0,
    parameter integer STATIC_PHASE3 = 0,
    parameter integer STATIC_PHASE4 = 0,
    parameter integer STATIC_PHASEPHY = 0,
    parameter integer STATIC_PHASEF = 0,
    parameter integer STATIC_CPHASE0 = 0,
    parameter integer STATIC_CPHASE1 = 0,
    parameter integer STATIC_CPHASE2 = 0,
    parameter integer STATIC_CPHASE3 = 0,
    parameter integer STATIC_CPHASE4 = 0,
    parameter integer STATIC_CPHASEPHY = 0,
    parameter integer STATIC_CPHASEF = 0,
    parameter CLKOUT0_SYN_EN = "FALSE",
    parameter CLKOUT1_SYN_EN = "FALSE",
    parameter CLKOUT2_SYN_EN = "FALSE",
    parameter CLKOUT3_SYN_EN = "FALSE",
    parameter CLKOUT4_SYN_EN = "FALSE",
    parameter CLKOUTPHY_SYN_EN = "FALSE",
    parameter CLKOUTF_SYN_EN = "FALSE",
    parameter INTERNAL_FB = "CLKOUTF",
    parameter EXTERNAL_FB = "DISABLE",
    parameter BANDWIDTH = "OPTIMIZED"
) (
    output CLKOUT0,
    output CLKOUT0N,
    output CLKOUT1,
    output CLKOUT1N,
    output CLKOUT2,
    output CLKOUT2N,
    output CLKOUT3,
    output CLKOUT3N,
    output CLKOUT4,
    output CLKOUTPHY,
    output CLKOUTPHYN,
    output CLKOUTF,
    output CLKOUTFN,
    output LOCK,
    output [15:0] APB_RDATA,
    output APB_READY,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUTPHY_SYN,
    input CLKOUTF_SYN,
    input PLL_PWD,
    input RST,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [15:0] APB_WDATA
)  ;
endmodule


module GTP_PPLL_DFT
#(
    parameter real CLKIN_FREQ = 50.0,
    parameter LOCK_MODE = 1'b0,
    parameter integer STATIC_RATIOI = 1,
    parameter integer STATIC_RATIOM = 1,
    parameter integer STATIC_RATIO0 = 1,
    parameter integer STATIC_RATIO1 = 1,
    parameter integer STATIC_RATIO2 = 1,
    parameter integer STATIC_RATIO3 = 1,
    parameter integer STATIC_RATIO4 = 1,
    parameter integer STATIC_RATIOPHY = 1,
    parameter integer STATIC_RATIOF = 1,
    parameter integer STATIC_DUTY0 = 2,
    parameter integer STATIC_DUTY1 = 2,
    parameter integer STATIC_DUTY2 = 2,
    parameter integer STATIC_DUTY3 = 2,
    parameter integer STATIC_DUTY4 = 2,
    parameter integer STATIC_DUTYPHY = 2,
    parameter integer STATIC_DUTYF = 2,
    parameter integer STATIC_PHASE0 = 0,
    parameter integer STATIC_PHASE1 = 0,
    parameter integer STATIC_PHASE2 = 0,
    parameter integer STATIC_PHASE3 = 0,
    parameter integer STATIC_PHASE4 = 0,
    parameter integer STATIC_PHASEPHY = 0,
    parameter integer STATIC_PHASEF = 0,
    parameter integer STATIC_CPHASE0 = 0,
    parameter integer STATIC_CPHASE1 = 0,
    parameter integer STATIC_CPHASE2 = 0,
    parameter integer STATIC_CPHASE3 = 0,
    parameter integer STATIC_CPHASE4 = 0,
    parameter integer STATIC_CPHASEPHY = 0,
    parameter integer STATIC_CPHASEF = 0,
    parameter CLKOUT0_SYN_EN = "FALSE",
    parameter CLKOUT1_SYN_EN = "FALSE",
    parameter CLKOUT2_SYN_EN = "FALSE",
    parameter CLKOUT3_SYN_EN = "FALSE",
    parameter CLKOUT4_SYN_EN = "FALSE",
    parameter CLKOUTPHY_SYN_EN = "FALSE",
    parameter CLKOUTF_SYN_EN = "FALSE",
    parameter INTERNAL_FB = "CLKOUTF",
    parameter EXTERNAL_FB = "DISABLE",
    parameter BANDWIDTH = "OPTIMIZED",
    parameter integer PFDTOP_CLKTEST_SEL = 0,
    parameter PFDTOP_CLKTEST_EN = "FALSE",
    parameter integer DCTEST_SEL = 0,
    parameter integer CP_CUR_SEL = 0,
    parameter VCTRL_TEST_EN = "FALSE"
) (
    output PFDTOP_CLK_TEST,
    output CLKOUT0,
    output CLKOUT0N,
    output CLKOUT1,
    output CLKOUT1N,
    output CLKOUT2,
    output CLKOUT2N,
    output CLKOUT3,
    output CLKOUT3N,
    output CLKOUT4,
    output CLKOUTPHY,
    output CLKOUTPHYN,
    output CLKOUTF,
    output CLKOUTFN,
    output LOCK,
    output [15:0] APB_RDATA,
    output APB_READY,
    input CLKIN1,
    input CLKIN2,
    input CLKFB,
    input CLKIN_SEL,
    input CLKOUT0_SYN,
    input CLKOUT1_SYN,
    input CLKOUT2_SYN,
    input CLKOUT3_SYN,
    input CLKOUT4_SYN,
    input CLKOUTPHY_SYN,
    input CLKOUTF_SYN,
    input PLL_PWD,
    input RST,
    input APB_CLK,
    input APB_RST_N,
    input [4:0] APB_ADDR,
    input APB_SEL,
    input APB_EN,
    input APB_WRITE,
    input [15:0] APB_WDATA
)  ;
endmodule


module GTP_RAM32X1DP
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output DO,
    input DI,
    input [4:0] RADDR,
    input [4:0] WADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM32X1SP
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output DO,
    input DI,
    input [4:0] ADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM32X2DP
#(
    parameter [31:0] INIT_0 = 32'h00000000,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] DO,
    input [1:0] DI,
    input [4:0] RADDR,
    input [4:0] WADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM32X2SP
#(
    parameter [31:0] INIT_0 = 32'h00000000,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] DO,
    input [1:0] DI,
    input [4:0] ADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM32X2X4
#(
    parameter [63:0] INIT_0 = 64'h0000000000000000,
    parameter [63:0] INIT_1 = 64'h0000000000000000,
    parameter [63:0] INIT_2 = 64'h0000000000000000,
    parameter [63:0] INIT_3 = 64'h0000000000000000
) (
    output [1:0] DO0,
    output [1:0] DO1,
    output [1:0] DO2,
    output [1:0] DO3,
    input [1:0] DI0,
    input [1:0] DI1,
    input [1:0] DI2,
    input [1:0] DI3,
    input [4:0] ADDR0,
    input [4:0] ADDR1,
    input [4:0] ADDR2,
    input [4:0] ADDR3,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM64X1DP
#(
    parameter [63:0] INIT = 64'h0000000000000000
) (
    output DO,
    input DI,
    input [5:0] RADDR,
    input [5:0] WADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM64X1SP
#(
    parameter [63:0] INIT = 64'h0000000000000000
) (
    output DO,
    input DI,
    input [5:0] ADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM64X1X4
#(
    parameter [63:0] INIT_0 = 64'h0000000000000000,
    parameter [63:0] INIT_1 = 64'h0000000000000000,
    parameter [63:0] INIT_2 = 64'h0000000000000000,
    parameter [63:0] INIT_3 = 64'h0000000000000000
) (
    output DO0,
    output DO1,
    output DO2,
    output DO3,
    input DI0,
    input DI1,
    input DI2,
    input DI3,
    input [5:0] ADDR0,
    input [5:0] ADDR1,
    input [5:0] ADDR2,
    input [5:0] ADDR3,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM128X1DP
#(
    parameter [127:0] INIT = 128'h00000000000000000000000000000000
) (
    output DO,
    input DI,
    input [6:0] RADDR,
    input [6:0] WADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM128X1SP
#(
    parameter [127:0] INIT = 128'h00000000000000000000000000000000
) (
    output DO,
    input DI,
    input [6:0] ADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RAM256X1SP
#(
    parameter [255:0] INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000
) (
    output DO,
    input DI,
    input [7:0] ADDR,
    input WCLK,
    input WE
)  ;
endmodule


module GTP_RES_CAL_E1
#(
    parameter CAL_ENABLE = "FALSE",
    parameter CAL_CASCADE = "LOCAL",
    parameter CASC_V_ENABLE = "FALSE",
    parameter BANK_LOC = "BANKR5"
) (
    input [4:0] PCODE_IN,
    input [4:0] NCODE_IN,
    input SAMPLE_IN,
    input EN,
    input CODE_SEL,
    input RST_N,
    output [4:0] PCODE_OUT,
    output [4:0] NCODE_OUT,
    output CAL_DONE
)  ;
endmodule


module GTP_RES_CAL_E1_DFT
#(
    parameter CAL_ENABLE = "FALSE",
    parameter CAL_CASCADE = "LOCAL",
    parameter CASC_V_ENABLE = "FALSE",
    parameter BANK_LOC = "BANKR5",
    parameter FAST_CAL_N = "FALSE"
) (
    input [4:0] PCODE_IN,
    input [4:0] NCODE_IN,
    input SAMPLE_IN,
    input EN,
    input CODE_SEL,
    input RST_N,
    output [4:0] PCODE_OUT,
    output [4:0] NCODE_OUT,
    output CAL_DONE
)  ;
endmodule


module GTP_RES_CAL_E2
#(
    parameter CAL_ENABLE = "FALSE",
    parameter CAL_CASCADE = "LOCAL",
    parameter CASC_V_ENABLE = "FALSE",
    parameter BANK_LOC = "BANKR5",
    parameter FAST_CAL_N = "FALSE"
) (
    input [4:0] PCODE_IN,
    input [4:0] NCODE_IN,
    input SAMPLE_IN,
    input EN,
    input CODE_SEL,
    input RST_N,
    output [4:0] PCODE_OUT,
    output [4:0] NCODE_OUT,
    output CAL_DONE
)  ;
endmodule


module GTP_ROM32X1
#(
    parameter [31:0] INIT = 32'h00000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4
)  ;
endmodule


module GTP_ROM32X2
#(
    parameter [31:0] INIT_0 = 32'h00000000,
    parameter [31:0] INIT_1 = 32'h00000000
) (
    output [1:0] Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4
)  ;
endmodule


module GTP_ROM64X1
#(
    parameter [63:0] INIT = 64'h0000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5
)  ;
endmodule


module GTP_ROM128X1
#(
    parameter [127:0] INIT = 128'h00000000000000000000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5,
    input I6
)  ;
endmodule


module GTP_ROM256X1
#(
    parameter [255:0] INIT = 256'h0000000000000000000000000000000000000000000000000000000000000000
) (
    output Z,
    input I0,
    input I1,
    input I2,
    input I3,
    input I4,
    input I5,
    input I6,
    input I7
)  ;
endmodule


module GTP_SCANCHAIN_E1
#(
    parameter [31:0] IDCODE = 32'hAAAA5555,
    parameter integer CHAIN_NUM = 1
) (
    output TDO,
    input TCK,
    input TDI,
    input TMS,
    output CAPDR,
    output SHFTDR,
    output UPDR,
    output JCLK,
    output RST,
    output JRTI,
    output FLG_USER,
    output TCK_USER,
    output TDI_USER,
    output TMS_USER,
    input TDO_USER
)  ;
endmodule


module GTP_START_E1
(
    output WAKEUP_OVER,
    input CLK,
    input GOE,
    input GRS_N,
    input GWE
)  ;
endmodule


module GTP_UDID
#(
    parameter integer UDID_WIDTH = 64,
    parameter [95:0] UDID_CODE = 96'h000000000000000000000000
) (
    input DI,
    output DO,
    input LOAD,
    input SE,
    input CLK
)  ;
endmodule


module GTP_ZERO
(
    output Z
)  ;
endmodule


module GTP_ZEROHOLDDELAY
#(
    parameter ZHOLD_SET = "NODELAY"
) (
    output DO,
    input DI
)  ;
endmodule

